module wallace_mult(a, b, prod_trim, exp);
input [31:0] a,b;
output [31:0] prod_trim;
wire [63:0] prod;
output exp;
wire a0b0, a0b1, a1b0, a0b2, a1b1, a2b0, a0b3, a1b2, a2b1, a3b0, a0b4, a1b3, a2b2, a3b1, a4b0, a0b5, a1b4, a2b3, a3b2, a4b1, a5b0, a0b6, a1b5, a2b4, a3b3, a4b2, a5b1, a6b0, a0b7, a1b6, a2b5, a3b4, a4b3, a5b2, a6b1, a7b0, a0b8, a1b7, a2b6, a3b5, a4b4, a5b3, a6b2, a7b1, a8b0, a0b9, a1b8, a2b7, a3b6, a4b5, a5b4, a6b3, a7b2, a8b1, a9b0, a0b10, a1b9, a2b8, a3b7, a4b6, a5b5, a6b4, a7b3, a8b2, a9b1, a10b0, a0b11, a1b10, a2b9, a3b8, a4b7, a5b6, a6b5, a7b4, a8b3, a9b2, a10b1, a11b0, a0b12, a1b11, a2b10, a3b9, a4b8, a5b7, a6b6, a7b5, a8b4, a9b3, a10b2, a11b1, a12b0, a0b13, a1b12, a2b11, a3b10, a4b9, a5b8, a6b7, a7b6, a8b5, a9b4, a10b3, a11b2, a12b1, a13b0, a0b14, a1b13, a2b12, a3b11, a4b10, a5b9, a6b8, a7b7, a8b6, a9b5, a10b4, a11b3, a12b2, a13b1, a14b0, a0b15, a1b14, a2b13, a3b12, a4b11, a5b10, a6b9, a7b8, a8b7, a9b6, a10b5, a11b4, a12b3, a13b2, a14b1, a15b0, a0b16, a1b15, a2b14, a3b13, a4b12, a5b11, a6b10, a7b9, a8b8, a9b7, a10b6, a11b5, a12b4, a13b3, a14b2, a15b1, a16b0, a0b17, a1b16, a2b15, a3b14, a4b13, a5b12, a6b11, a7b10, a8b9, a9b8, a10b7, a11b6, a12b5, a13b4, a14b3, a15b2, a16b1, a17b0, a0b18, a1b17, a2b16, a3b15, a4b14, a5b13, a6b12, a7b11, a8b10, a9b9, a10b8, a11b7, a12b6, a13b5, a14b4, a15b3, a16b2, a17b1, a18b0, a0b19, a1b18, a2b17, a3b16, a4b15, a5b14, a6b13, a7b12, a8b11, a9b10, a10b9, a11b8, a12b7, a13b6, a14b5, a15b4, a16b3, a17b2, a18b1, a19b0, a0b20, a1b19, a2b18, a3b17, a4b16, a5b15, a6b14, a7b13, a8b12, a9b11, a10b10, a11b9, a12b8, a13b7, a14b6, a15b5, a16b4, a17b3, a18b2, a19b1, a20b0, a0b21, a1b20, a2b19, a3b18, a4b17, a5b16, a6b15, a7b14, a8b13, a9b12, a10b11, a11b10, a12b9, a13b8, a14b7, a15b6, a16b5, a17b4, a18b3, a19b2, a20b1, a21b0, a0b22, a1b21, a2b20, a3b19, a4b18, a5b17, a6b16, a7b15, a8b14, a9b13, a10b12, a11b11, a12b10, a13b9, a14b8, a15b7, a16b6, a17b5, a18b4, a19b3, a20b2, a21b1, a22b0, a0b23, a1b22, a2b21, a3b20, a4b19, a5b18, a6b17, a7b16, a8b15, a9b14, a10b13, a11b12, a12b11, a13b10, a14b9, a15b8, a16b7, a17b6, a18b5, a19b4, a20b3, a21b2, a22b1, a23b0, a0b24, a1b23, a2b22, a3b21, a4b20, a5b19, a6b18, a7b17, a8b16, a9b15, a10b14, a11b13, a12b12, a13b11, a14b10, a15b9, a16b8, a17b7, a18b6, a19b5, a20b4, a21b3, a22b2, a23b1, a24b0, a0b25, a1b24, a2b23, a3b22, a4b21, a5b20, a6b19, a7b18, a8b17, a9b16, a10b15, a11b14, a12b13, a13b12, a14b11, a15b10, a16b9, a17b8, a18b7, a19b6, a20b5, a21b4, a22b3, a23b2, a24b1, a25b0, a0b26, a1b25, a2b24, a3b23, a4b22, a5b21, a6b20, a7b19, a8b18, a9b17, a10b16, a11b15, a12b14, a13b13, a14b12, a15b11, a16b10, a17b9, a18b8, a19b7, a20b6, a21b5, a22b4, a23b3, a24b2, a25b1, a26b0, a0b27, a1b26, a2b25, a3b24, a4b23, a5b22, a6b21, a7b20, a8b19, a9b18, a10b17, a11b16, a12b15, a13b14, a14b13, a15b12, a16b11, a17b10, a18b9, a19b8, a20b7, a21b6, a22b5, a23b4, a24b3, a25b2, a26b1, a27b0, a0b28, a1b27, a2b26, a3b25, a4b24, a5b23, a6b22, a7b21, a8b20, a9b19, a10b18, a11b17, a12b16, a13b15, a14b14, a15b13, a16b12, a17b11, a18b10, a19b9, a20b8, a21b7, a22b6, a23b5, a24b4, a25b3, a26b2, a27b1, a28b0, a0b29, a1b28, a2b27, a3b26, a4b25, a5b24, a6b23, a7b22, a8b21, a9b20, a10b19, a11b18, a12b17, a13b16, a14b15, a15b14, a16b13, a17b12, a18b11, a19b10, a20b9, a21b8, a22b7, a23b6, a24b5, a25b4, a26b3, a27b2, a28b1, a29b0, a0b30, a1b29, a2b28, a3b27, a4b26, a5b25, a6b24, a7b23, a8b22, a9b21, a10b20, a11b19, a12b18, a13b17, a14b16, a15b15, a16b14, a17b13, a18b12, a19b11, a20b10, a21b9, a22b8, a23b7, a24b6, a25b5, a26b4, a27b3, a28b2, a29b1, a30b0, a0b31, a1b30, a2b29, a3b28, a4b27, a5b26, a6b25, a7b24, a8b23, a9b22, a10b21, a11b20, a12b19, a13b18, a14b17, a15b16, a16b15, a17b14, a18b13, a19b12, a20b11, a21b10, a22b9, a23b8, a24b7, a25b6, a26b5, a27b4, a28b3, a29b2, a30b1, a31b0;

//Weight 1
assign a0b0 = a[0]&b[0];

//Weight 2
assign a0b1 = a[0]&b[1];
assign a1b0 = a[1]&b[0];

//Weight 4
assign a0b2 = a[0]&b[2];
assign a1b1 = a[1]&b[1];
assign a2b0 = a[2]&b[0];

//Weight 8
assign a0b3 = a[0]&b[3];
assign a1b2 = a[1]&b[2];
assign a2b1 = a[2]&b[1];
assign a3b0 = a[3]&b[0];

//Weight 16
assign a0b4 = a[0]&b[4];
assign a1b3 = a[1]&b[3];
assign a2b2 = a[2]&b[2];
assign a3b1 = a[3]&b[1];
assign a4b0 = a[4]&b[0];

//Weight 32
assign a0b5 = a[0]&b[5];
assign a1b4 = a[1]&b[4];
assign a2b3 = a[2]&b[3];
assign a3b2 = a[3]&b[2];
assign a4b1 = a[4]&b[1];
assign a5b0 = a[5]&b[0];

//Weight 64
assign a0b6 = a[0]&b[6];
assign a1b5 = a[1]&b[5];
assign a2b4 = a[2]&b[4];
assign a3b3 = a[3]&b[3];
assign a4b2 = a[4]&b[2];
assign a5b1 = a[5]&b[1];
assign a6b0 = a[6]&b[0];

//Weight 128
assign a0b7 = a[0]&b[7];
assign a1b6 = a[1]&b[6];
assign a2b5 = a[2]&b[5];
assign a3b4 = a[3]&b[4];
assign a4b3 = a[4]&b[3];
assign a5b2 = a[5]&b[2];
assign a6b1 = a[6]&b[1];
assign a7b0 = a[7]&b[0];

//Weight 256
assign a0b8 = a[0]&b[8];
assign a1b7 = a[1]&b[7];
assign a2b6 = a[2]&b[6];
assign a3b5 = a[3]&b[5];
assign a4b4 = a[4]&b[4];
assign a5b3 = a[5]&b[3];
assign a6b2 = a[6]&b[2];
assign a7b1 = a[7]&b[1];
assign a8b0 = a[8]&b[0];

//Weight 512
assign a0b9 = a[0]&b[9];
assign a1b8 = a[1]&b[8];
assign a2b7 = a[2]&b[7];
assign a3b6 = a[3]&b[6];
assign a4b5 = a[4]&b[5];
assign a5b4 = a[5]&b[4];
assign a6b3 = a[6]&b[3];
assign a7b2 = a[7]&b[2];
assign a8b1 = a[8]&b[1];
assign a9b0 = a[9]&b[0];

//Weight 1024
assign a0b10 = a[0]&b[10];
assign a1b9 = a[1]&b[9];
assign a2b8 = a[2]&b[8];
assign a3b7 = a[3]&b[7];
assign a4b6 = a[4]&b[6];
assign a5b5 = a[5]&b[5];
assign a6b4 = a[6]&b[4];
assign a7b3 = a[7]&b[3];
assign a8b2 = a[8]&b[2];
assign a9b1 = a[9]&b[1];
assign a10b0 = a[10]&b[0];

//Weight 2048
assign a0b11 = a[0]&b[11];
assign a1b10 = a[1]&b[10];
assign a2b9 = a[2]&b[9];
assign a3b8 = a[3]&b[8];
assign a4b7 = a[4]&b[7];
assign a5b6 = a[5]&b[6];
assign a6b5 = a[6]&b[5];
assign a7b4 = a[7]&b[4];
assign a8b3 = a[8]&b[3];
assign a9b2 = a[9]&b[2];
assign a10b1 = a[10]&b[1];
assign a11b0 = a[11]&b[0];

//Weight 4096
assign a0b12 = a[0]&b[12];
assign a1b11 = a[1]&b[11];
assign a2b10 = a[2]&b[10];
assign a3b9 = a[3]&b[9];
assign a4b8 = a[4]&b[8];
assign a5b7 = a[5]&b[7];
assign a6b6 = a[6]&b[6];
assign a7b5 = a[7]&b[5];
assign a8b4 = a[8]&b[4];
assign a9b3 = a[9]&b[3];
assign a10b2 = a[10]&b[2];
assign a11b1 = a[11]&b[1];
assign a12b0 = a[12]&b[0];

//Weight 8192
assign a0b13 = a[0]&b[13];
assign a1b12 = a[1]&b[12];
assign a2b11 = a[2]&b[11];
assign a3b10 = a[3]&b[10];
assign a4b9 = a[4]&b[9];
assign a5b8 = a[5]&b[8];
assign a6b7 = a[6]&b[7];
assign a7b6 = a[7]&b[6];
assign a8b5 = a[8]&b[5];
assign a9b4 = a[9]&b[4];
assign a10b3 = a[10]&b[3];
assign a11b2 = a[11]&b[2];
assign a12b1 = a[12]&b[1];
assign a13b0 = a[13]&b[0];

//Weight 16384
assign a0b14 = a[0]&b[14];
assign a1b13 = a[1]&b[13];
assign a2b12 = a[2]&b[12];
assign a3b11 = a[3]&b[11];
assign a4b10 = a[4]&b[10];
assign a5b9 = a[5]&b[9];
assign a6b8 = a[6]&b[8];
assign a7b7 = a[7]&b[7];
assign a8b6 = a[8]&b[6];
assign a9b5 = a[9]&b[5];
assign a10b4 = a[10]&b[4];
assign a11b3 = a[11]&b[3];
assign a12b2 = a[12]&b[2];
assign a13b1 = a[13]&b[1];
assign a14b0 = a[14]&b[0];

//Weight 32768
assign a0b15 = a[0]&b[15];
assign a1b14 = a[1]&b[14];
assign a2b13 = a[2]&b[13];
assign a3b12 = a[3]&b[12];
assign a4b11 = a[4]&b[11];
assign a5b10 = a[5]&b[10];
assign a6b9 = a[6]&b[9];
assign a7b8 = a[7]&b[8];
assign a8b7 = a[8]&b[7];
assign a9b6 = a[9]&b[6];
assign a10b5 = a[10]&b[5];
assign a11b4 = a[11]&b[4];
assign a12b3 = a[12]&b[3];
assign a13b2 = a[13]&b[2];
assign a14b1 = a[14]&b[1];
assign a15b0 = a[15]&b[0];

//Weight 65536
assign a0b16 = a[0]&b[16];
assign a1b15 = a[1]&b[15];
assign a2b14 = a[2]&b[14];
assign a3b13 = a[3]&b[13];
assign a4b12 = a[4]&b[12];
assign a5b11 = a[5]&b[11];
assign a6b10 = a[6]&b[10];
assign a7b9 = a[7]&b[9];
assign a8b8 = a[8]&b[8];
assign a9b7 = a[9]&b[7];
assign a10b6 = a[10]&b[6];
assign a11b5 = a[11]&b[5];
assign a12b4 = a[12]&b[4];
assign a13b3 = a[13]&b[3];
assign a14b2 = a[14]&b[2];
assign a15b1 = a[15]&b[1];
assign a16b0 = a[16]&b[0];

//Weight 131072
assign a0b17 = a[0]&b[17];
assign a1b16 = a[1]&b[16];
assign a2b15 = a[2]&b[15];
assign a3b14 = a[3]&b[14];
assign a4b13 = a[4]&b[13];
assign a5b12 = a[5]&b[12];
assign a6b11 = a[6]&b[11];
assign a7b10 = a[7]&b[10];
assign a8b9 = a[8]&b[9];
assign a9b8 = a[9]&b[8];
assign a10b7 = a[10]&b[7];
assign a11b6 = a[11]&b[6];
assign a12b5 = a[12]&b[5];
assign a13b4 = a[13]&b[4];
assign a14b3 = a[14]&b[3];
assign a15b2 = a[15]&b[2];
assign a16b1 = a[16]&b[1];
assign a17b0 = a[17]&b[0];

//Weight 262144
assign a0b18 = a[0]&b[18];
assign a1b17 = a[1]&b[17];
assign a2b16 = a[2]&b[16];
assign a3b15 = a[3]&b[15];
assign a4b14 = a[4]&b[14];
assign a5b13 = a[5]&b[13];
assign a6b12 = a[6]&b[12];
assign a7b11 = a[7]&b[11];
assign a8b10 = a[8]&b[10];
assign a9b9 = a[9]&b[9];
assign a10b8 = a[10]&b[8];
assign a11b7 = a[11]&b[7];
assign a12b6 = a[12]&b[6];
assign a13b5 = a[13]&b[5];
assign a14b4 = a[14]&b[4];
assign a15b3 = a[15]&b[3];
assign a16b2 = a[16]&b[2];
assign a17b1 = a[17]&b[1];
assign a18b0 = a[18]&b[0];

//Weight 524288
assign a0b19 = a[0]&b[19];
assign a1b18 = a[1]&b[18];
assign a2b17 = a[2]&b[17];
assign a3b16 = a[3]&b[16];
assign a4b15 = a[4]&b[15];
assign a5b14 = a[5]&b[14];
assign a6b13 = a[6]&b[13];
assign a7b12 = a[7]&b[12];
assign a8b11 = a[8]&b[11];
assign a9b10 = a[9]&b[10];
assign a10b9 = a[10]&b[9];
assign a11b8 = a[11]&b[8];
assign a12b7 = a[12]&b[7];
assign a13b6 = a[13]&b[6];
assign a14b5 = a[14]&b[5];
assign a15b4 = a[15]&b[4];
assign a16b3 = a[16]&b[3];
assign a17b2 = a[17]&b[2];
assign a18b1 = a[18]&b[1];
assign a19b0 = a[19]&b[0];

//Weight 1048576
assign a0b20 = a[0]&b[20];
assign a1b19 = a[1]&b[19];
assign a2b18 = a[2]&b[18];
assign a3b17 = a[3]&b[17];
assign a4b16 = a[4]&b[16];
assign a5b15 = a[5]&b[15];
assign a6b14 = a[6]&b[14];
assign a7b13 = a[7]&b[13];
assign a8b12 = a[8]&b[12];
assign a9b11 = a[9]&b[11];
assign a10b10 = a[10]&b[10];
assign a11b9 = a[11]&b[9];
assign a12b8 = a[12]&b[8];
assign a13b7 = a[13]&b[7];
assign a14b6 = a[14]&b[6];
assign a15b5 = a[15]&b[5];
assign a16b4 = a[16]&b[4];
assign a17b3 = a[17]&b[3];
assign a18b2 = a[18]&b[2];
assign a19b1 = a[19]&b[1];
assign a20b0 = a[20]&b[0];

//Weight 2097152
assign a0b21 = a[0]&b[21];
assign a1b20 = a[1]&b[20];
assign a2b19 = a[2]&b[19];
assign a3b18 = a[3]&b[18];
assign a4b17 = a[4]&b[17];
assign a5b16 = a[5]&b[16];
assign a6b15 = a[6]&b[15];
assign a7b14 = a[7]&b[14];
assign a8b13 = a[8]&b[13];
assign a9b12 = a[9]&b[12];
assign a10b11 = a[10]&b[11];
assign a11b10 = a[11]&b[10];
assign a12b9 = a[12]&b[9];
assign a13b8 = a[13]&b[8];
assign a14b7 = a[14]&b[7];
assign a15b6 = a[15]&b[6];
assign a16b5 = a[16]&b[5];
assign a17b4 = a[17]&b[4];
assign a18b3 = a[18]&b[3];
assign a19b2 = a[19]&b[2];
assign a20b1 = a[20]&b[1];
assign a21b0 = a[21]&b[0];

//Weight 4194304
assign a0b22 = a[0]&b[22];
assign a1b21 = a[1]&b[21];
assign a2b20 = a[2]&b[20];
assign a3b19 = a[3]&b[19];
assign a4b18 = a[4]&b[18];
assign a5b17 = a[5]&b[17];
assign a6b16 = a[6]&b[16];
assign a7b15 = a[7]&b[15];
assign a8b14 = a[8]&b[14];
assign a9b13 = a[9]&b[13];
assign a10b12 = a[10]&b[12];
assign a11b11 = a[11]&b[11];
assign a12b10 = a[12]&b[10];
assign a13b9 = a[13]&b[9];
assign a14b8 = a[14]&b[8];
assign a15b7 = a[15]&b[7];
assign a16b6 = a[16]&b[6];
assign a17b5 = a[17]&b[5];
assign a18b4 = a[18]&b[4];
assign a19b3 = a[19]&b[3];
assign a20b2 = a[20]&b[2];
assign a21b1 = a[21]&b[1];
assign a22b0 = a[22]&b[0];

//Weight 8388608
assign a0b23 = a[0]&b[23];
assign a1b22 = a[1]&b[22];
assign a2b21 = a[2]&b[21];
assign a3b20 = a[3]&b[20];
assign a4b19 = a[4]&b[19];
assign a5b18 = a[5]&b[18];
assign a6b17 = a[6]&b[17];
assign a7b16 = a[7]&b[16];
assign a8b15 = a[8]&b[15];
assign a9b14 = a[9]&b[14];
assign a10b13 = a[10]&b[13];
assign a11b12 = a[11]&b[12];
assign a12b11 = a[12]&b[11];
assign a13b10 = a[13]&b[10];
assign a14b9 = a[14]&b[9];
assign a15b8 = a[15]&b[8];
assign a16b7 = a[16]&b[7];
assign a17b6 = a[17]&b[6];
assign a18b5 = a[18]&b[5];
assign a19b4 = a[19]&b[4];
assign a20b3 = a[20]&b[3];
assign a21b2 = a[21]&b[2];
assign a22b1 = a[22]&b[1];
assign a23b0 = a[23]&b[0];

//Weight 16777216
assign a0b24 = a[0]&b[24];
assign a1b23 = a[1]&b[23];
assign a2b22 = a[2]&b[22];
assign a3b21 = a[3]&b[21];
assign a4b20 = a[4]&b[20];
assign a5b19 = a[5]&b[19];
assign a6b18 = a[6]&b[18];
assign a7b17 = a[7]&b[17];
assign a8b16 = a[8]&b[16];
assign a9b15 = a[9]&b[15];
assign a10b14 = a[10]&b[14];
assign a11b13 = a[11]&b[13];
assign a12b12 = a[12]&b[12];
assign a13b11 = a[13]&b[11];
assign a14b10 = a[14]&b[10];
assign a15b9 = a[15]&b[9];
assign a16b8 = a[16]&b[8];
assign a17b7 = a[17]&b[7];
assign a18b6 = a[18]&b[6];
assign a19b5 = a[19]&b[5];
assign a20b4 = a[20]&b[4];
assign a21b3 = a[21]&b[3];
assign a22b2 = a[22]&b[2];
assign a23b1 = a[23]&b[1];
assign a24b0 = a[24]&b[0];

//Weight 33554432
assign a0b25 = a[0]&b[25];
assign a1b24 = a[1]&b[24];
assign a2b23 = a[2]&b[23];
assign a3b22 = a[3]&b[22];
assign a4b21 = a[4]&b[21];
assign a5b20 = a[5]&b[20];
assign a6b19 = a[6]&b[19];
assign a7b18 = a[7]&b[18];
assign a8b17 = a[8]&b[17];
assign a9b16 = a[9]&b[16];
assign a10b15 = a[10]&b[15];
assign a11b14 = a[11]&b[14];
assign a12b13 = a[12]&b[13];
assign a13b12 = a[13]&b[12];
assign a14b11 = a[14]&b[11];
assign a15b10 = a[15]&b[10];
assign a16b9 = a[16]&b[9];
assign a17b8 = a[17]&b[8];
assign a18b7 = a[18]&b[7];
assign a19b6 = a[19]&b[6];
assign a20b5 = a[20]&b[5];
assign a21b4 = a[21]&b[4];
assign a22b3 = a[22]&b[3];
assign a23b2 = a[23]&b[2];
assign a24b1 = a[24]&b[1];
assign a25b0 = a[25]&b[0];

//Weight 67108864
assign a0b26 = a[0]&b[26];
assign a1b25 = a[1]&b[25];
assign a2b24 = a[2]&b[24];
assign a3b23 = a[3]&b[23];
assign a4b22 = a[4]&b[22];
assign a5b21 = a[5]&b[21];
assign a6b20 = a[6]&b[20];
assign a7b19 = a[7]&b[19];
assign a8b18 = a[8]&b[18];
assign a9b17 = a[9]&b[17];
assign a10b16 = a[10]&b[16];
assign a11b15 = a[11]&b[15];
assign a12b14 = a[12]&b[14];
assign a13b13 = a[13]&b[13];
assign a14b12 = a[14]&b[12];
assign a15b11 = a[15]&b[11];
assign a16b10 = a[16]&b[10];
assign a17b9 = a[17]&b[9];
assign a18b8 = a[18]&b[8];
assign a19b7 = a[19]&b[7];
assign a20b6 = a[20]&b[6];
assign a21b5 = a[21]&b[5];
assign a22b4 = a[22]&b[4];
assign a23b3 = a[23]&b[3];
assign a24b2 = a[24]&b[2];
assign a25b1 = a[25]&b[1];
assign a26b0 = a[26]&b[0];

//Weight 134217728
assign a0b27 = a[0]&b[27];
assign a1b26 = a[1]&b[26];
assign a2b25 = a[2]&b[25];
assign a3b24 = a[3]&b[24];
assign a4b23 = a[4]&b[23];
assign a5b22 = a[5]&b[22];
assign a6b21 = a[6]&b[21];
assign a7b20 = a[7]&b[20];
assign a8b19 = a[8]&b[19];
assign a9b18 = a[9]&b[18];
assign a10b17 = a[10]&b[17];
assign a11b16 = a[11]&b[16];
assign a12b15 = a[12]&b[15];
assign a13b14 = a[13]&b[14];
assign a14b13 = a[14]&b[13];
assign a15b12 = a[15]&b[12];
assign a16b11 = a[16]&b[11];
assign a17b10 = a[17]&b[10];
assign a18b9 = a[18]&b[9];
assign a19b8 = a[19]&b[8];
assign a20b7 = a[20]&b[7];
assign a21b6 = a[21]&b[6];
assign a22b5 = a[22]&b[5];
assign a23b4 = a[23]&b[4];
assign a24b3 = a[24]&b[3];
assign a25b2 = a[25]&b[2];
assign a26b1 = a[26]&b[1];
assign a27b0 = a[27]&b[0];

//Weight 268435456
assign a0b28 = a[0]&b[28];
assign a1b27 = a[1]&b[27];
assign a2b26 = a[2]&b[26];
assign a3b25 = a[3]&b[25];
assign a4b24 = a[4]&b[24];
assign a5b23 = a[5]&b[23];
assign a6b22 = a[6]&b[22];
assign a7b21 = a[7]&b[21];
assign a8b20 = a[8]&b[20];
assign a9b19 = a[9]&b[19];
assign a10b18 = a[10]&b[18];
assign a11b17 = a[11]&b[17];
assign a12b16 = a[12]&b[16];
assign a13b15 = a[13]&b[15];
assign a14b14 = a[14]&b[14];
assign a15b13 = a[15]&b[13];
assign a16b12 = a[16]&b[12];
assign a17b11 = a[17]&b[11];
assign a18b10 = a[18]&b[10];
assign a19b9 = a[19]&b[9];
assign a20b8 = a[20]&b[8];
assign a21b7 = a[21]&b[7];
assign a22b6 = a[22]&b[6];
assign a23b5 = a[23]&b[5];
assign a24b4 = a[24]&b[4];
assign a25b3 = a[25]&b[3];
assign a26b2 = a[26]&b[2];
assign a27b1 = a[27]&b[1];
assign a28b0 = a[28]&b[0];

//Weight 536870912
assign a0b29 = a[0]&b[29];
assign a1b28 = a[1]&b[28];
assign a2b27 = a[2]&b[27];
assign a3b26 = a[3]&b[26];
assign a4b25 = a[4]&b[25];
assign a5b24 = a[5]&b[24];
assign a6b23 = a[6]&b[23];
assign a7b22 = a[7]&b[22];
assign a8b21 = a[8]&b[21];
assign a9b20 = a[9]&b[20];
assign a10b19 = a[10]&b[19];
assign a11b18 = a[11]&b[18];
assign a12b17 = a[12]&b[17];
assign a13b16 = a[13]&b[16];
assign a14b15 = a[14]&b[15];
assign a15b14 = a[15]&b[14];
assign a16b13 = a[16]&b[13];
assign a17b12 = a[17]&b[12];
assign a18b11 = a[18]&b[11];
assign a19b10 = a[19]&b[10];
assign a20b9 = a[20]&b[9];
assign a21b8 = a[21]&b[8];
assign a22b7 = a[22]&b[7];
assign a23b6 = a[23]&b[6];
assign a24b5 = a[24]&b[5];
assign a25b4 = a[25]&b[4];
assign a26b3 = a[26]&b[3];
assign a27b2 = a[27]&b[2];
assign a28b1 = a[28]&b[1];
assign a29b0 = a[29]&b[0];

//Weight 1073741824
assign a0b30 = a[0]&b[30];
assign a1b29 = a[1]&b[29];
assign a2b28 = a[2]&b[28];
assign a3b27 = a[3]&b[27];
assign a4b26 = a[4]&b[26];
assign a5b25 = a[5]&b[25];
assign a6b24 = a[6]&b[24];
assign a7b23 = a[7]&b[23];
assign a8b22 = a[8]&b[22];
assign a9b21 = a[9]&b[21];
assign a10b20 = a[10]&b[20];
assign a11b19 = a[11]&b[19];
assign a12b18 = a[12]&b[18];
assign a13b17 = a[13]&b[17];
assign a14b16 = a[14]&b[16];
assign a15b15 = a[15]&b[15];
assign a16b14 = a[16]&b[14];
assign a17b13 = a[17]&b[13];
assign a18b12 = a[18]&b[12];
assign a19b11 = a[19]&b[11];
assign a20b10 = a[20]&b[10];
assign a21b9 = a[21]&b[9];
assign a22b8 = a[22]&b[8];
assign a23b7 = a[23]&b[7];
assign a24b6 = a[24]&b[6];
assign a25b5 = a[25]&b[5];
assign a26b4 = a[26]&b[4];
assign a27b3 = a[27]&b[3];
assign a28b2 = a[28]&b[2];
assign a29b1 = a[29]&b[1];
assign a30b0 = a[30]&b[0];

//Weight 2147483648
assign a0b31 = ~(a[0]&b[31]);
assign a1b30 = a[1]&b[30];
assign a2b29 = a[2]&b[29];
assign a3b28 = a[3]&b[28];
assign a4b27 = a[4]&b[27];
assign a5b26 = a[5]&b[26];
assign a6b25 = a[6]&b[25];
assign a7b24 = a[7]&b[24];
assign a8b23 = a[8]&b[23];
assign a9b22 = a[9]&b[22];
assign a10b21 = a[10]&b[21];
assign a11b20 = a[11]&b[20];
assign a12b19 = a[12]&b[19];
assign a13b18 = a[13]&b[18];
assign a14b17 = a[14]&b[17];
assign a15b16 = a[15]&b[16];
assign a16b15 = a[16]&b[15];
assign a17b14 = a[17]&b[14];
assign a18b13 = a[18]&b[13];
assign a19b12 = a[19]&b[12];
assign a20b11 = a[20]&b[11];
assign a21b10 = a[21]&b[10];
assign a22b9 = a[22]&b[9];
assign a23b8 = a[23]&b[8];
assign a24b7 = a[24]&b[7];
assign a25b6 = a[25]&b[6];
assign a26b5 = a[26]&b[5];
assign a27b4 = a[27]&b[4];
assign a28b3 = a[28]&b[3];
assign a29b2 = a[29]&b[2];
assign a30b1 = a[30]&b[1];
assign a31b0 = ~(a[31]&b[0]);

//Weight 4294967296
assign a1b31 = ~(a[1]&b[31]);
assign a2b30 = a[2]&b[30];
assign a3b29 = a[3]&b[29];
assign a4b28 = a[4]&b[28];
assign a5b27 = a[5]&b[27];
assign a6b26 = a[6]&b[26];
assign a7b25 = a[7]&b[25];
assign a8b24 = a[8]&b[24];
assign a9b23 = a[9]&b[23];
assign a10b22 = a[10]&b[22];
assign a11b21 = a[11]&b[21];
assign a12b20 = a[12]&b[20];
assign a13b19 = a[13]&b[19];
assign a14b18 = a[14]&b[18];
assign a15b17 = a[15]&b[17];
assign a16b16 = a[16]&b[16];
assign a17b15 = a[17]&b[15];
assign a18b14 = a[18]&b[14];
assign a19b13 = a[19]&b[13];
assign a20b12 = a[20]&b[12];
assign a21b11 = a[21]&b[11];
assign a22b10 = a[22]&b[10];
assign a23b9 = a[23]&b[9];
assign a24b8 = a[24]&b[8];
assign a25b7 = a[25]&b[7];
assign a26b6 = a[26]&b[6];
assign a27b5 = a[27]&b[5];
assign a28b4 = a[28]&b[4];
assign a29b3 = a[29]&b[3];
assign a30b2 = a[30]&b[2];
assign a31b1 = ~(a[31]&b[1]);

//Weight 8589934592
assign a2b31 = ~(a[2]&b[31]);
assign a3b30 = a[3]&b[30];
assign a4b29 = a[4]&b[29];
assign a5b28 = a[5]&b[28];
assign a6b27 = a[6]&b[27];
assign a7b26 = a[7]&b[26];
assign a8b25 = a[8]&b[25];
assign a9b24 = a[9]&b[24];
assign a10b23 = a[10]&b[23];
assign a11b22 = a[11]&b[22];
assign a12b21 = a[12]&b[21];
assign a13b20 = a[13]&b[20];
assign a14b19 = a[14]&b[19];
assign a15b18 = a[15]&b[18];
assign a16b17 = a[16]&b[17];
assign a17b16 = a[17]&b[16];
assign a18b15 = a[18]&b[15];
assign a19b14 = a[19]&b[14];
assign a20b13 = a[20]&b[13];
assign a21b12 = a[21]&b[12];
assign a22b11 = a[22]&b[11];
assign a23b10 = a[23]&b[10];
assign a24b9 = a[24]&b[9];
assign a25b8 = a[25]&b[8];
assign a26b7 = a[26]&b[7];
assign a27b6 = a[27]&b[6];
assign a28b5 = a[28]&b[5];
assign a29b4 = a[29]&b[4];
assign a30b3 = a[30]&b[3];
assign a31b2 = ~(a[31]&b[2]);

//Weight 17179869184
assign a3b31 = ~(a[3]&b[31]);
assign a4b30 = a[4]&b[30];
assign a5b29 = a[5]&b[29];
assign a6b28 = a[6]&b[28];
assign a7b27 = a[7]&b[27];
assign a8b26 = a[8]&b[26];
assign a9b25 = a[9]&b[25];
assign a10b24 = a[10]&b[24];
assign a11b23 = a[11]&b[23];
assign a12b22 = a[12]&b[22];
assign a13b21 = a[13]&b[21];
assign a14b20 = a[14]&b[20];
assign a15b19 = a[15]&b[19];
assign a16b18 = a[16]&b[18];
assign a17b17 = a[17]&b[17];
assign a18b16 = a[18]&b[16];
assign a19b15 = a[19]&b[15];
assign a20b14 = a[20]&b[14];
assign a21b13 = a[21]&b[13];
assign a22b12 = a[22]&b[12];
assign a23b11 = a[23]&b[11];
assign a24b10 = a[24]&b[10];
assign a25b9 = a[25]&b[9];
assign a26b8 = a[26]&b[8];
assign a27b7 = a[27]&b[7];
assign a28b6 = a[28]&b[6];
assign a29b5 = a[29]&b[5];
assign a30b4 = a[30]&b[4];
assign a31b3 = ~(a[31]&b[3]);

//Weight 34359738368
assign a4b31 = ~(a[4]&b[31]);
assign a5b30 = a[5]&b[30];
assign a6b29 = a[6]&b[29];
assign a7b28 = a[7]&b[28];
assign a8b27 = a[8]&b[27];
assign a9b26 = a[9]&b[26];
assign a10b25 = a[10]&b[25];
assign a11b24 = a[11]&b[24];
assign a12b23 = a[12]&b[23];
assign a13b22 = a[13]&b[22];
assign a14b21 = a[14]&b[21];
assign a15b20 = a[15]&b[20];
assign a16b19 = a[16]&b[19];
assign a17b18 = a[17]&b[18];
assign a18b17 = a[18]&b[17];
assign a19b16 = a[19]&b[16];
assign a20b15 = a[20]&b[15];
assign a21b14 = a[21]&b[14];
assign a22b13 = a[22]&b[13];
assign a23b12 = a[23]&b[12];
assign a24b11 = a[24]&b[11];
assign a25b10 = a[25]&b[10];
assign a26b9 = a[26]&b[9];
assign a27b8 = a[27]&b[8];
assign a28b7 = a[28]&b[7];
assign a29b6 = a[29]&b[6];
assign a30b5 = a[30]&b[5];
assign a31b4 = ~(a[31]&b[4]);

//Weight 68719476736
assign a5b31 = ~(a[5]&b[31]);
assign a6b30 = a[6]&b[30];
assign a7b29 = a[7]&b[29];
assign a8b28 = a[8]&b[28];
assign a9b27 = a[9]&b[27];
assign a10b26 = a[10]&b[26];
assign a11b25 = a[11]&b[25];
assign a12b24 = a[12]&b[24];
assign a13b23 = a[13]&b[23];
assign a14b22 = a[14]&b[22];
assign a15b21 = a[15]&b[21];
assign a16b20 = a[16]&b[20];
assign a17b19 = a[17]&b[19];
assign a18b18 = a[18]&b[18];
assign a19b17 = a[19]&b[17];
assign a20b16 = a[20]&b[16];
assign a21b15 = a[21]&b[15];
assign a22b14 = a[22]&b[14];
assign a23b13 = a[23]&b[13];
assign a24b12 = a[24]&b[12];
assign a25b11 = a[25]&b[11];
assign a26b10 = a[26]&b[10];
assign a27b9 = a[27]&b[9];
assign a28b8 = a[28]&b[8];
assign a29b7 = a[29]&b[7];
assign a30b6 = a[30]&b[6];
assign a31b5 = ~(a[31]&b[5]);

//Weight 137438953472
assign a6b31 = ~(a[6]&b[31]);
assign a7b30 = a[7]&b[30];
assign a8b29 = a[8]&b[29];
assign a9b28 = a[9]&b[28];
assign a10b27 = a[10]&b[27];
assign a11b26 = a[11]&b[26];
assign a12b25 = a[12]&b[25];
assign a13b24 = a[13]&b[24];
assign a14b23 = a[14]&b[23];
assign a15b22 = a[15]&b[22];
assign a16b21 = a[16]&b[21];
assign a17b20 = a[17]&b[20];
assign a18b19 = a[18]&b[19];
assign a19b18 = a[19]&b[18];
assign a20b17 = a[20]&b[17];
assign a21b16 = a[21]&b[16];
assign a22b15 = a[22]&b[15];
assign a23b14 = a[23]&b[14];
assign a24b13 = a[24]&b[13];
assign a25b12 = a[25]&b[12];
assign a26b11 = a[26]&b[11];
assign a27b10 = a[27]&b[10];
assign a28b9 = a[28]&b[9];
assign a29b8 = a[29]&b[8];
assign a30b7 = a[30]&b[7];
assign a31b6 = ~(a[31]&b[6]);

//Weight 274877906944
assign a7b31 = ~(a[7]&b[31]);
assign a8b30 = a[8]&b[30];
assign a9b29 = a[9]&b[29];
assign a10b28 = a[10]&b[28];
assign a11b27 = a[11]&b[27];
assign a12b26 = a[12]&b[26];
assign a13b25 = a[13]&b[25];
assign a14b24 = a[14]&b[24];
assign a15b23 = a[15]&b[23];
assign a16b22 = a[16]&b[22];
assign a17b21 = a[17]&b[21];
assign a18b20 = a[18]&b[20];
assign a19b19 = a[19]&b[19];
assign a20b18 = a[20]&b[18];
assign a21b17 = a[21]&b[17];
assign a22b16 = a[22]&b[16];
assign a23b15 = a[23]&b[15];
assign a24b14 = a[24]&b[14];
assign a25b13 = a[25]&b[13];
assign a26b12 = a[26]&b[12];
assign a27b11 = a[27]&b[11];
assign a28b10 = a[28]&b[10];
assign a29b9 = a[29]&b[9];
assign a30b8 = a[30]&b[8];
assign a31b7 = ~(a[31]&b[7]);

//Weight 549755813888
assign a8b31 = ~(a[8]&b[31]);
assign a9b30 = a[9]&b[30];
assign a10b29 = a[10]&b[29];
assign a11b28 = a[11]&b[28];
assign a12b27 = a[12]&b[27];
assign a13b26 = a[13]&b[26];
assign a14b25 = a[14]&b[25];
assign a15b24 = a[15]&b[24];
assign a16b23 = a[16]&b[23];
assign a17b22 = a[17]&b[22];
assign a18b21 = a[18]&b[21];
assign a19b20 = a[19]&b[20];
assign a20b19 = a[20]&b[19];
assign a21b18 = a[21]&b[18];
assign a22b17 = a[22]&b[17];
assign a23b16 = a[23]&b[16];
assign a24b15 = a[24]&b[15];
assign a25b14 = a[25]&b[14];
assign a26b13 = a[26]&b[13];
assign a27b12 = a[27]&b[12];
assign a28b11 = a[28]&b[11];
assign a29b10 = a[29]&b[10];
assign a30b9 = a[30]&b[9];
assign a31b8 = ~(a[31]&b[8]);

//Weight 1099511627776
assign a9b31 = ~(a[9]&b[31]);
assign a10b30 = a[10]&b[30];
assign a11b29 = a[11]&b[29];
assign a12b28 = a[12]&b[28];
assign a13b27 = a[13]&b[27];
assign a14b26 = a[14]&b[26];
assign a15b25 = a[15]&b[25];
assign a16b24 = a[16]&b[24];
assign a17b23 = a[17]&b[23];
assign a18b22 = a[18]&b[22];
assign a19b21 = a[19]&b[21];
assign a20b20 = a[20]&b[20];
assign a21b19 = a[21]&b[19];
assign a22b18 = a[22]&b[18];
assign a23b17 = a[23]&b[17];
assign a24b16 = a[24]&b[16];
assign a25b15 = a[25]&b[15];
assign a26b14 = a[26]&b[14];
assign a27b13 = a[27]&b[13];
assign a28b12 = a[28]&b[12];
assign a29b11 = a[29]&b[11];
assign a30b10 = a[30]&b[10];
assign a31b9 = ~(a[31]&b[9]);

//Weight 2199023255552
assign a10b31 = ~(a[10]&b[31]);
assign a11b30 = a[11]&b[30];
assign a12b29 = a[12]&b[29];
assign a13b28 = a[13]&b[28];
assign a14b27 = a[14]&b[27];
assign a15b26 = a[15]&b[26];
assign a16b25 = a[16]&b[25];
assign a17b24 = a[17]&b[24];
assign a18b23 = a[18]&b[23];
assign a19b22 = a[19]&b[22];
assign a20b21 = a[20]&b[21];
assign a21b20 = a[21]&b[20];
assign a22b19 = a[22]&b[19];
assign a23b18 = a[23]&b[18];
assign a24b17 = a[24]&b[17];
assign a25b16 = a[25]&b[16];
assign a26b15 = a[26]&b[15];
assign a27b14 = a[27]&b[14];
assign a28b13 = a[28]&b[13];
assign a29b12 = a[29]&b[12];
assign a30b11 = a[30]&b[11];
assign a31b10 = ~(a[31]&b[10]);

//Weight 4398046511104
assign a11b31 = ~(a[11]&b[31]);
assign a12b30 = a[12]&b[30];
assign a13b29 = a[13]&b[29];
assign a14b28 = a[14]&b[28];
assign a15b27 = a[15]&b[27];
assign a16b26 = a[16]&b[26];
assign a17b25 = a[17]&b[25];
assign a18b24 = a[18]&b[24];
assign a19b23 = a[19]&b[23];
assign a20b22 = a[20]&b[22];
assign a21b21 = a[21]&b[21];
assign a22b20 = a[22]&b[20];
assign a23b19 = a[23]&b[19];
assign a24b18 = a[24]&b[18];
assign a25b17 = a[25]&b[17];
assign a26b16 = a[26]&b[16];
assign a27b15 = a[27]&b[15];
assign a28b14 = a[28]&b[14];
assign a29b13 = a[29]&b[13];
assign a30b12 = a[30]&b[12];
assign a31b11 = ~(a[31]&b[11]);

//Weight 8796093022208
assign a12b31 = ~(a[12]&b[31]);
assign a13b30 = a[13]&b[30];
assign a14b29 = a[14]&b[29];
assign a15b28 = a[15]&b[28];
assign a16b27 = a[16]&b[27];
assign a17b26 = a[17]&b[26];
assign a18b25 = a[18]&b[25];
assign a19b24 = a[19]&b[24];
assign a20b23 = a[20]&b[23];
assign a21b22 = a[21]&b[22];
assign a22b21 = a[22]&b[21];
assign a23b20 = a[23]&b[20];
assign a24b19 = a[24]&b[19];
assign a25b18 = a[25]&b[18];
assign a26b17 = a[26]&b[17];
assign a27b16 = a[27]&b[16];
assign a28b15 = a[28]&b[15];
assign a29b14 = a[29]&b[14];
assign a30b13 = a[30]&b[13];
assign a31b12 = ~(a[31]&b[12]);

//Weight 17592186044416
assign a13b31 = ~(a[13]&b[31]);
assign a14b30 = a[14]&b[30];
assign a15b29 = a[15]&b[29];
assign a16b28 = a[16]&b[28];
assign a17b27 = a[17]&b[27];
assign a18b26 = a[18]&b[26];
assign a19b25 = a[19]&b[25];
assign a20b24 = a[20]&b[24];
assign a21b23 = a[21]&b[23];
assign a22b22 = a[22]&b[22];
assign a23b21 = a[23]&b[21];
assign a24b20 = a[24]&b[20];
assign a25b19 = a[25]&b[19];
assign a26b18 = a[26]&b[18];
assign a27b17 = a[27]&b[17];
assign a28b16 = a[28]&b[16];
assign a29b15 = a[29]&b[15];
assign a30b14 = a[30]&b[14];
assign a31b13 = ~(a[31]&b[13]);

//Weight 35184372088832
assign a14b31 = ~(a[14]&b[31]);
assign a15b30 = a[15]&b[30];
assign a16b29 = a[16]&b[29];
assign a17b28 = a[17]&b[28];
assign a18b27 = a[18]&b[27];
assign a19b26 = a[19]&b[26];
assign a20b25 = a[20]&b[25];
assign a21b24 = a[21]&b[24];
assign a22b23 = a[22]&b[23];
assign a23b22 = a[23]&b[22];
assign a24b21 = a[24]&b[21];
assign a25b20 = a[25]&b[20];
assign a26b19 = a[26]&b[19];
assign a27b18 = a[27]&b[18];
assign a28b17 = a[28]&b[17];
assign a29b16 = a[29]&b[16];
assign a30b15 = a[30]&b[15];
assign a31b14 = ~(a[31]&b[14]);

//Weight 70368744177664
assign a15b31 = ~(a[15]&b[31]);
assign a16b30 = a[16]&b[30];
assign a17b29 = a[17]&b[29];
assign a18b28 = a[18]&b[28];
assign a19b27 = a[19]&b[27];
assign a20b26 = a[20]&b[26];
assign a21b25 = a[21]&b[25];
assign a22b24 = a[22]&b[24];
assign a23b23 = a[23]&b[23];
assign a24b22 = a[24]&b[22];
assign a25b21 = a[25]&b[21];
assign a26b20 = a[26]&b[20];
assign a27b19 = a[27]&b[19];
assign a28b18 = a[28]&b[18];
assign a29b17 = a[29]&b[17];
assign a30b16 = a[30]&b[16];
assign a31b15 = ~(a[31]&b[15]);

//Weight 140737488355328
assign a16b31 = ~(a[16]&b[31]);
assign a17b30 = a[17]&b[30];
assign a18b29 = a[18]&b[29];
assign a19b28 = a[19]&b[28];
assign a20b27 = a[20]&b[27];
assign a21b26 = a[21]&b[26];
assign a22b25 = a[22]&b[25];
assign a23b24 = a[23]&b[24];
assign a24b23 = a[24]&b[23];
assign a25b22 = a[25]&b[22];
assign a26b21 = a[26]&b[21];
assign a27b20 = a[27]&b[20];
assign a28b19 = a[28]&b[19];
assign a29b18 = a[29]&b[18];
assign a30b17 = a[30]&b[17];
assign a31b16 = ~(a[31]&b[16]);

//Weight 281474976710656
assign a17b31 = ~(a[17]&b[31]);
assign a18b30 = a[18]&b[30];
assign a19b29 = a[19]&b[29];
assign a20b28 = a[20]&b[28];
assign a21b27 = a[21]&b[27];
assign a22b26 = a[22]&b[26];
assign a23b25 = a[23]&b[25];
assign a24b24 = a[24]&b[24];
assign a25b23 = a[25]&b[23];
assign a26b22 = a[26]&b[22];
assign a27b21 = a[27]&b[21];
assign a28b20 = a[28]&b[20];
assign a29b19 = a[29]&b[19];
assign a30b18 = a[30]&b[18];
assign a31b17 = ~(a[31]&b[17]);

//Weight 562949953421312
assign a18b31 = ~(a[18]&b[31]);
assign a19b30 = a[19]&b[30];
assign a20b29 = a[20]&b[29];
assign a21b28 = a[21]&b[28];
assign a22b27 = a[22]&b[27];
assign a23b26 = a[23]&b[26];
assign a24b25 = a[24]&b[25];
assign a25b24 = a[25]&b[24];
assign a26b23 = a[26]&b[23];
assign a27b22 = a[27]&b[22];
assign a28b21 = a[28]&b[21];
assign a29b20 = a[29]&b[20];
assign a30b19 = a[30]&b[19];
assign a31b18 = ~(a[31]&b[18]);

//Weight 1125899906842624
assign a19b31 = ~(a[19]&b[31]);
assign a20b30 = a[20]&b[30];
assign a21b29 = a[21]&b[29];
assign a22b28 = a[22]&b[28];
assign a23b27 = a[23]&b[27];
assign a24b26 = a[24]&b[26];
assign a25b25 = a[25]&b[25];
assign a26b24 = a[26]&b[24];
assign a27b23 = a[27]&b[23];
assign a28b22 = a[28]&b[22];
assign a29b21 = a[29]&b[21];
assign a30b20 = a[30]&b[20];
assign a31b19 = ~(a[31]&b[19]);

//Weight 2251799813685248
assign a20b31 = ~(a[20]&b[31]);
assign a21b30 = a[21]&b[30];
assign a22b29 = a[22]&b[29];
assign a23b28 = a[23]&b[28];
assign a24b27 = a[24]&b[27];
assign a25b26 = a[25]&b[26];
assign a26b25 = a[26]&b[25];
assign a27b24 = a[27]&b[24];
assign a28b23 = a[28]&b[23];
assign a29b22 = a[29]&b[22];
assign a30b21 = a[30]&b[21];
assign a31b20 = ~(a[31]&b[20]);

//Weight 4503599627370496
assign a21b31 = ~(a[21]&b[31]);
assign a22b30 = a[22]&b[30];
assign a23b29 = a[23]&b[29];
assign a24b28 = a[24]&b[28];
assign a25b27 = a[25]&b[27];
assign a26b26 = a[26]&b[26];
assign a27b25 = a[27]&b[25];
assign a28b24 = a[28]&b[24];
assign a29b23 = a[29]&b[23];
assign a30b22 = a[30]&b[22];
assign a31b21 = ~(a[31]&b[21]);

//Weight 9007199254740992
assign a22b31 = ~(a[22]&b[31]);
assign a23b30 = a[23]&b[30];
assign a24b29 = a[24]&b[29];
assign a25b28 = a[25]&b[28];
assign a26b27 = a[26]&b[27];
assign a27b26 = a[27]&b[26];
assign a28b25 = a[28]&b[25];
assign a29b24 = a[29]&b[24];
assign a30b23 = a[30]&b[23];
assign a31b22 = ~(a[31]&b[22]);

//Weight 18014398509481984
assign a23b31 = ~(a[23]&b[31]);
assign a24b30 = a[24]&b[30];
assign a25b29 = a[25]&b[29];
assign a26b28 = a[26]&b[28];
assign a27b27 = a[27]&b[27];
assign a28b26 = a[28]&b[26];
assign a29b25 = a[29]&b[25];
assign a30b24 = a[30]&b[24];
assign a31b23 = ~(a[31]&b[23]);

//Weight 36028797018963968
assign a24b31 = ~(a[24]&b[31]);
assign a25b30 = a[25]&b[30];
assign a26b29 = a[26]&b[29];
assign a27b28 = a[27]&b[28];
assign a28b27 = a[28]&b[27];
assign a29b26 = a[29]&b[26];
assign a30b25 = a[30]&b[25];
assign a31b24 = ~(a[31]&b[24]);

//Weight 72057594037927936
assign a25b31 = ~(a[25]&b[31]);
assign a26b30 = a[26]&b[30];
assign a27b29 = a[27]&b[29];
assign a28b28 = a[28]&b[28];
assign a29b27 = a[29]&b[27];
assign a30b26 = a[30]&b[26];
assign a31b25 = ~(a[31]&b[25]);

//Weight 144115188075855872
assign a26b31 = ~(a[26]&b[31]);
assign a27b30 = a[27]&b[30];
assign a28b29 = a[28]&b[29];
assign a29b28 = a[29]&b[28];
assign a30b27 = a[30]&b[27];
assign a31b26 = ~(a[31]&b[26]);

//Weight 288230376151711744
assign a27b31 = ~(a[27]&b[31]);
assign a28b30 = a[28]&b[30];
assign a29b29 = a[29]&b[29];
assign a30b28 = a[30]&b[28];
assign a31b27 = ~(a[31]&b[27]);

//Weight 576460752303423488
assign a28b31 = ~(a[28]&b[31]);
assign a29b30 = a[29]&b[30];
assign a30b29 = a[30]&b[29];
assign a31b28 = ~(a[31]&b[28]);

//Weight 1152921504606846976
assign a29b31 = ~(a[29]&b[31]);
assign a30b30 = a[30]&b[30];
assign a31b29 = ~(a[31]&b[29]);

//Weight 2305843009213693952
assign a30b31 = ~(a[30]&b[31]);
assign a31b30 = ~(a[31]&b[30]);

//Weight 4611686018427387904
assign a31b31 = (a[31]&b[31]);

//Weight 9223372036854775808

//[['a0b0'], ['a0b1', 'a1b0'], ['a0b2', 'a1b1', 'a2b0'], ['a0b3', 'a1b2', 'a2b1', 'a3b0'], ['a0b4', 'a1b3', 'a2b2', 'a3b1', 'a4b0'], ['a0b5', 'a1b4', 'a2b3', 'a3b2', 'a4b1', 'a5b0'], ['a0b6', 'a1b5', 'a2b4', 'a3b3', 'a4b2', 'a5b1', 'a6b0'], ['a0b7', 'a1b6', 'a2b5', 'a3b4', 'a4b3', 'a5b2', 'a6b1', 'a7b0'], ['a0b8', 'a1b7', 'a2b6', 'a3b5', 'a4b4', 'a5b3', 'a6b2', 'a7b1', 'a8b0'], ['a0b9', 'a1b8', 'a2b7', 'a3b6', 'a4b5', 'a5b4', 'a6b3', 'a7b2', 'a8b1', 'a9b0'], ['a0b10', 'a1b9', 'a2b8', 'a3b7', 'a4b6', 'a5b5', 'a6b4', 'a7b3', 'a8b2', 'a9b1', 'a10b0'], ['a0b11', 'a1b10', 'a2b9', 'a3b8', 'a4b7', 'a5b6', 'a6b5', 'a7b4', 'a8b3', 'a9b2', 'a10b1', 'a11b0'], ['a0b12', 'a1b11', 'a2b10', 'a3b9', 'a4b8', 'a5b7', 'a6b6', 'a7b5', 'a8b4', 'a9b3', 'a10b2', 'a11b1', 'a12b0'], ['a0b13', 'a1b12', 'a2b11', 'a3b10', 'a4b9', 'a5b8', 'a6b7', 'a7b6', 'a8b5', 'a9b4', 'a10b3', 'a11b2', 'a12b1', 'a13b0'], ['a0b14', 'a1b13', 'a2b12', 'a3b11', 'a4b10', 'a5b9', 'a6b8', 'a7b7', 'a8b6', 'a9b5', 'a10b4', 'a11b3', 'a12b2', 'a13b1', 'a14b0'], ['a0b15', 'a1b14', 'a2b13', 'a3b12', 'a4b11', 'a5b10', 'a6b9', 'a7b8', 'a8b7', 'a9b6', 'a10b5', 'a11b4', 'a12b3', 'a13b2', 'a14b1', 'a15b0'], ['a0b16', 'a1b15', 'a2b14', 'a3b13', 'a4b12', 'a5b11', 'a6b10', 'a7b9', 'a8b8', 'a9b7', 'a10b6', 'a11b5', 'a12b4', 'a13b3', 'a14b2', 'a15b1', 'a16b0'], ['a0b17', 'a1b16', 'a2b15', 'a3b14', 'a4b13', 'a5b12', 'a6b11', 'a7b10', 'a8b9', 'a9b8', 'a10b7', 'a11b6', 'a12b5', 'a13b4', 'a14b3', 'a15b2', 'a16b1', 'a17b0'], ['a0b18', 'a1b17', 'a2b16', 'a3b15', 'a4b14', 'a5b13', 'a6b12', 'a7b11', 'a8b10', 'a9b9', 'a10b8', 'a11b7', 'a12b6', 'a13b5', 'a14b4', 'a15b3', 'a16b2', 'a17b1', 'a18b0'], ['a0b19', 'a1b18', 'a2b17', 'a3b16', 'a4b15', 'a5b14', 'a6b13', 'a7b12', 'a8b11', 'a9b10', 'a10b9', 'a11b8', 'a12b7', 'a13b6', 'a14b5', 'a15b4', 'a16b3', 'a17b2', 'a18b1', 'a19b0'], ['a0b20', 'a1b19', 'a2b18', 'a3b17', 'a4b16', 'a5b15', 'a6b14', 'a7b13', 'a8b12', 'a9b11', 'a10b10', 'a11b9', 'a12b8', 'a13b7', 'a14b6', 'a15b5', 'a16b4', 'a17b3', 'a18b2', 'a19b1', 'a20b0'], ['a0b21', 'a1b20', 'a2b19', 'a3b18', 'a4b17', 'a5b16', 'a6b15', 'a7b14', 'a8b13', 'a9b12', 'a10b11', 'a11b10', 'a12b9', 'a13b8', 'a14b7', 'a15b6', 'a16b5', 'a17b4', 'a18b3', 'a19b2', 'a20b1', 'a21b0'], ['a0b22', 'a1b21', 'a2b20', 'a3b19', 'a4b18', 'a5b17', 'a6b16', 'a7b15', 'a8b14', 'a9b13', 'a10b12', 'a11b11', 'a12b10', 'a13b9', 'a14b8', 'a15b7', 'a16b6', 'a17b5', 'a18b4', 'a19b3', 'a20b2', 'a21b1', 'a22b0'], ['a0b23', 'a1b22', 'a2b21', 'a3b20', 'a4b19', 'a5b18', 'a6b17', 'a7b16', 'a8b15', 'a9b14', 'a10b13', 'a11b12', 'a12b11', 'a13b10', 'a14b9', 'a15b8', 'a16b7', 'a17b6', 'a18b5', 'a19b4', 'a20b3', 'a21b2', 'a22b1', 'a23b0'], ['a0b24', 'a1b23', 'a2b22', 'a3b21', 'a4b20', 'a5b19', 'a6b18', 'a7b17', 'a8b16', 'a9b15', 'a10b14', 'a11b13', 'a12b12', 'a13b11', 'a14b10', 'a15b9', 'a16b8', 'a17b7', 'a18b6', 'a19b5', 'a20b4', 'a21b3', 'a22b2', 'a23b1', 'a24b0'], ['a0b25', 'a1b24', 'a2b23', 'a3b22', 'a4b21', 'a5b20', 'a6b19', 'a7b18', 'a8b17', 'a9b16', 'a10b15', 'a11b14', 'a12b13', 'a13b12', 'a14b11', 'a15b10', 'a16b9', 'a17b8', 'a18b7', 'a19b6', 'a20b5', 'a21b4', 'a22b3', 'a23b2', 'a24b1', 'a25b0'], ['a0b26', 'a1b25', 'a2b24', 'a3b23', 'a4b22', 'a5b21', 'a6b20', 'a7b19', 'a8b18', 'a9b17', 'a10b16', 'a11b15', 'a12b14', 'a13b13', 'a14b12', 'a15b11', 'a16b10', 'a17b9', 'a18b8', 'a19b7', 'a20b6', 'a21b5', 'a22b4', 'a23b3', 'a24b2', 'a25b1', 'a26b0'], ['a0b27', 'a1b26', 'a2b25', 'a3b24', 'a4b23', 'a5b22', 'a6b21', 'a7b20', 'a8b19', 'a9b18', 'a10b17', 'a11b16', 'a12b15', 'a13b14', 'a14b13', 'a15b12', 'a16b11', 'a17b10', 'a18b9', 'a19b8', 'a20b7', 'a21b6', 'a22b5', 'a23b4', 'a24b3', 'a25b2', 'a26b1', 'a27b0'], ['a0b28', 'a1b27', 'a2b26', 'a3b25', 'a4b24', 'a5b23', 'a6b22', 'a7b21', 'a8b20', 'a9b19', 'a10b18', 'a11b17', 'a12b16', 'a13b15', 'a14b14', 'a15b13', 'a16b12', 'a17b11', 'a18b10', 'a19b9', 'a20b8', 'a21b7', 'a22b6', 'a23b5', 'a24b4', 'a25b3', 'a26b2', 'a27b1', 'a28b0'], ['a0b29', 'a1b28', 'a2b27', 'a3b26', 'a4b25', 'a5b24', 'a6b23', 'a7b22', 'a8b21', 'a9b20', 'a10b19', 'a11b18', 'a12b17', 'a13b16', 'a14b15', 'a15b14', 'a16b13', 'a17b12', 'a18b11', 'a19b10', 'a20b9', 'a21b8', 'a22b7', 'a23b6', 'a24b5', 'a25b4', 'a26b3', 'a27b2', 'a28b1', 'a29b0'], ['a0b30', 'a1b29', 'a2b28', 'a3b27', 'a4b26', 'a5b25', 'a6b24', 'a7b23', 'a8b22', 'a9b21', 'a10b20', 'a11b19', 'a12b18', 'a13b17', 'a14b16', 'a15b15', 'a16b14', 'a17b13', 'a18b12', 'a19b11', 'a20b10', 'a21b9', 'a22b8', 'a23b7', 'a24b6', 'a25b5', 'a26b4', 'a27b3', 'a28b2', 'a29b1', 'a30b0'], ['a0b31', 'a1b30', 'a2b29', 'a3b28', 'a4b27', 'a5b26', 'a6b25', 'a7b24', 'a8b23', 'a9b22', 'a10b21', 'a11b20', 'a12b19', 'a13b18', 'a14b17', 'a15b16', 'a16b15', 'a17b14', 'a18b13', 'a19b12', 'a20b11', 'a21b10', 'a22b9', 'a23b8', 'a24b7', 'a25b6', 'a26b5', 'a27b4', 'a28b3', 'a29b2', 'a30b1', 'a31b0'], ['a1b31', 'a2b30', 'a3b29', 'a4b28', 'a5b27', 'a6b26', 'a7b25', 'a8b24', 'a9b23', 'a10b22', 'a11b21', 'a12b20', 'a13b19', 'a14b18', 'a15b17', 'a16b16', 'a17b15', 'a18b14', 'a19b13', 'a20b12', 'a21b11', 'a22b10', 'a23b9', 'a24b8', 'a25b7', 'a26b6', 'a27b5', 'a28b4', 'a29b3', 'a30b2', 'a31b1', "1'b1"], ['a2b31', 'a3b30', 'a4b29', 'a5b28', 'a6b27', 'a7b26', 'a8b25', 'a9b24', 'a10b23', 'a11b22', 'a12b21', 'a13b20', 'a14b19', 'a15b18', 'a16b17', 'a17b16', 'a18b15', 'a19b14', 'a20b13', 'a21b12', 'a22b11', 'a23b10', 'a24b9', 'a25b8', 'a26b7', 'a27b6', 'a28b5', 'a29b4', 'a30b3', 'a31b2'], ['a3b31', 'a4b30', 'a5b29', 'a6b28', 'a7b27', 'a8b26', 'a9b25', 'a10b24', 'a11b23', 'a12b22', 'a13b21', 'a14b20', 'a15b19', 'a16b18', 'a17b17', 'a18b16', 'a19b15', 'a20b14', 'a21b13', 'a22b12', 'a23b11', 'a24b10', 'a25b9', 'a26b8', 'a27b7', 'a28b6', 'a29b5', 'a30b4', 'a31b3'], ['a4b31', 'a5b30', 'a6b29', 'a7b28', 'a8b27', 'a9b26', 'a10b25', 'a11b24', 'a12b23', 'a13b22', 'a14b21', 'a15b20', 'a16b19', 'a17b18', 'a18b17', 'a19b16', 'a20b15', 'a21b14', 'a22b13', 'a23b12', 'a24b11', 'a25b10', 'a26b9', 'a27b8', 'a28b7', 'a29b6', 'a30b5', 'a31b4'], ['a5b31', 'a6b30', 'a7b29', 'a8b28', 'a9b27', 'a10b26', 'a11b25', 'a12b24', 'a13b23', 'a14b22', 'a15b21', 'a16b20', 'a17b19', 'a18b18', 'a19b17', 'a20b16', 'a21b15', 'a22b14', 'a23b13', 'a24b12', 'a25b11', 'a26b10', 'a27b9', 'a28b8', 'a29b7', 'a30b6', 'a31b5'], ['a6b31', 'a7b30', 'a8b29', 'a9b28', 'a10b27', 'a11b26', 'a12b25', 'a13b24', 'a14b23', 'a15b22', 'a16b21', 'a17b20', 'a18b19', 'a19b18', 'a20b17', 'a21b16', 'a22b15', 'a23b14', 'a24b13', 'a25b12', 'a26b11', 'a27b10', 'a28b9', 'a29b8', 'a30b7', 'a31b6'], ['a7b31', 'a8b30', 'a9b29', 'a10b28', 'a11b27', 'a12b26', 'a13b25', 'a14b24', 'a15b23', 'a16b22', 'a17b21', 'a18b20', 'a19b19', 'a20b18', 'a21b17', 'a22b16', 'a23b15', 'a24b14', 'a25b13', 'a26b12', 'a27b11', 'a28b10', 'a29b9', 'a30b8', 'a31b7'], ['a8b31', 'a9b30', 'a10b29', 'a11b28', 'a12b27', 'a13b26', 'a14b25', 'a15b24', 'a16b23', 'a17b22', 'a18b21', 'a19b20', 'a20b19', 'a21b18', 'a22b17', 'a23b16', 'a24b15', 'a25b14', 'a26b13', 'a27b12', 'a28b11', 'a29b10', 'a30b9', 'a31b8'], ['a9b31', 'a10b30', 'a11b29', 'a12b28', 'a13b27', 'a14b26', 'a15b25', 'a16b24', 'a17b23', 'a18b22', 'a19b21', 'a20b20', 'a21b19', 'a22b18', 'a23b17', 'a24b16', 'a25b15', 'a26b14', 'a27b13', 'a28b12', 'a29b11', 'a30b10', 'a31b9'], ['a10b31', 'a11b30', 'a12b29', 'a13b28', 'a14b27', 'a15b26', 'a16b25', 'a17b24', 'a18b23', 'a19b22', 'a20b21', 'a21b20', 'a22b19', 'a23b18', 'a24b17', 'a25b16', 'a26b15', 'a27b14', 'a28b13', 'a29b12', 'a30b11', 'a31b10'], ['a11b31', 'a12b30', 'a13b29', 'a14b28', 'a15b27', 'a16b26', 'a17b25', 'a18b24', 'a19b23', 'a20b22', 'a21b21', 'a22b20', 'a23b19', 'a24b18', 'a25b17', 'a26b16', 'a27b15', 'a28b14', 'a29b13', 'a30b12', 'a31b11'], ['a12b31', 'a13b30', 'a14b29', 'a15b28', 'a16b27', 'a17b26', 'a18b25', 'a19b24', 'a20b23', 'a21b22', 'a22b21', 'a23b20', 'a24b19', 'a25b18', 'a26b17', 'a27b16', 'a28b15', 'a29b14', 'a30b13', 'a31b12'], ['a13b31', 'a14b30', 'a15b29', 'a16b28', 'a17b27', 'a18b26', 'a19b25', 'a20b24', 'a21b23', 'a22b22', 'a23b21', 'a24b20', 'a25b19', 'a26b18', 'a27b17', 'a28b16', 'a29b15', 'a30b14', 'a31b13'], ['a14b31', 'a15b30', 'a16b29', 'a17b28', 'a18b27', 'a19b26', 'a20b25', 'a21b24', 'a22b23', 'a23b22', 'a24b21', 'a25b20', 'a26b19', 'a27b18', 'a28b17', 'a29b16', 'a30b15', 'a31b14'], ['a15b31', 'a16b30', 'a17b29', 'a18b28', 'a19b27', 'a20b26', 'a21b25', 'a22b24', 'a23b23', 'a24b22', 'a25b21', 'a26b20', 'a27b19', 'a28b18', 'a29b17', 'a30b16', 'a31b15'], ['a16b31', 'a17b30', 'a18b29', 'a19b28', 'a20b27', 'a21b26', 'a22b25', 'a23b24', 'a24b23', 'a25b22', 'a26b21', 'a27b20', 'a28b19', 'a29b18', 'a30b17', 'a31b16'], ['a17b31', 'a18b30', 'a19b29', 'a20b28', 'a21b27', 'a22b26', 'a23b25', 'a24b24', 'a25b23', 'a26b22', 'a27b21', 'a28b20', 'a29b19', 'a30b18', 'a31b17'], ['a18b31', 'a19b30', 'a20b29', 'a21b28', 'a22b27', 'a23b26', 'a24b25', 'a25b24', 'a26b23', 'a27b22', 'a28b21', 'a29b20', 'a30b19', 'a31b18'], ['a19b31', 'a20b30', 'a21b29', 'a22b28', 'a23b27', 'a24b26', 'a25b25', 'a26b24', 'a27b23', 'a28b22', 'a29b21', 'a30b20', 'a31b19'], ['a20b31', 'a21b30', 'a22b29', 'a23b28', 'a24b27', 'a25b26', 'a26b25', 'a27b24', 'a28b23', 'a29b22', 'a30b21', 'a31b20'], ['a21b31', 'a22b30', 'a23b29', 'a24b28', 'a25b27', 'a26b26', 'a27b25', 'a28b24', 'a29b23', 'a30b22', 'a31b21'], ['a22b31', 'a23b30', 'a24b29', 'a25b28', 'a26b27', 'a27b26', 'a28b25', 'a29b24', 'a30b23', 'a31b22'], ['a23b31', 'a24b30', 'a25b29', 'a26b28', 'a27b27', 'a28b26', 'a29b25', 'a30b24', 'a31b23'], ['a24b31', 'a25b30', 'a26b29', 'a27b28', 'a28b27', 'a29b26', 'a30b25', 'a31b24'], ['a25b31', 'a26b30', 'a27b29', 'a28b28', 'a29b27', 'a30b26', 'a31b25'], ['a26b31', 'a27b30', 'a28b29', 'a29b28', 'a30b27', 'a31b26'], ['a27b31', 'a28b30', 'a29b29', 'a30b28', 'a31b27'], ['a28b31', 'a29b30', 'a30b29', 'a31b28'], ['a29b31', 'a30b30', 'a31b29'], ['a30b31', 'a31b30'], ['a31b31'], ["1'b1"]]
assign prod[0] = a0b0;

wire lay1_ha0_s, lay1_ha0_c;
half_adder lay1_ha0(a1b0, a0b1, lay1_ha0_s, lay1_ha0_c);
assign prod[1] = lay1_ha0_s;

wire lay2_fa0_s, lay2_fa0_c;
full_adder lay2_fa0(a2b0, a1b1, a0b2, lay2_fa0_s, lay2_fa0_c);
wire lay2_ha0_s, lay2_ha0_c;
half_adder lay2_ha0(lay2_fa0_s, lay1_ha0_c, lay2_ha0_s, lay2_ha0_c);
assign prod[2] = lay2_ha0_s;

wire lay3_fa0_s, lay3_fa0_c;
full_adder lay3_fa0(a3b0, a2b1, a1b2, lay3_fa0_s, lay3_fa0_c);
wire lay3_fa1_s, lay3_fa1_c;
full_adder lay3_fa1(lay3_fa0_s, a0b3, lay2_ha0_c, lay3_fa1_s, lay3_fa1_c);
wire lay3_ha0_s, lay3_ha0_c;
half_adder lay3_ha0(lay3_fa1_s, lay2_fa0_c, lay3_ha0_s, lay3_ha0_c);
assign prod[3] = lay3_ha0_s;

wire lay4_fa0_s, lay4_fa0_c;
full_adder lay4_fa0(a4b0, a3b1, a2b2, lay4_fa0_s, lay4_fa0_c);
wire lay4_fa1_s, lay4_fa1_c;
full_adder lay4_fa1(lay4_fa0_s, a1b3, a0b4, lay4_fa1_s, lay4_fa1_c);
wire lay4_fa2_s, lay4_fa2_c;
full_adder lay4_fa2(lay4_fa1_s, lay3_ha0_c, lay3_fa1_c, lay4_fa2_s, lay4_fa2_c);
wire lay4_ha0_s, lay4_ha0_c;
half_adder lay4_ha0(lay4_fa2_s, lay3_fa0_c, lay4_ha0_s, lay4_ha0_c);
assign prod[4] = lay4_ha0_s;

wire lay5_fa0_s, lay5_fa0_c;
full_adder lay5_fa0(a5b0, a4b1, a3b2, lay5_fa0_s, lay5_fa0_c);
wire lay5_fa1_s, lay5_fa1_c;
full_adder lay5_fa1(lay5_fa0_s, a2b3, a1b4, lay5_fa1_s, lay5_fa1_c);
wire lay5_fa2_s, lay5_fa2_c;
full_adder lay5_fa2(lay5_fa1_s, a0b5, lay4_ha0_c, lay5_fa2_s, lay5_fa2_c);
wire lay5_fa3_s, lay5_fa3_c;
full_adder lay5_fa3(lay5_fa2_s, lay4_fa2_c, lay4_fa1_c, lay5_fa3_s, lay5_fa3_c);
wire lay5_ha0_s, lay5_ha0_c;
half_adder lay5_ha0(lay5_fa3_s, lay4_fa0_c, lay5_ha0_s, lay5_ha0_c);
assign prod[5] = lay5_ha0_s;

wire lay6_fa0_s, lay6_fa0_c;
full_adder lay6_fa0(a6b0, a5b1, a4b2, lay6_fa0_s, lay6_fa0_c);
wire lay6_fa1_s, lay6_fa1_c;
full_adder lay6_fa1(lay6_fa0_s, a3b3, a2b4, lay6_fa1_s, lay6_fa1_c);
wire lay6_fa2_s, lay6_fa2_c;
full_adder lay6_fa2(lay6_fa1_s, a1b5, a0b6, lay6_fa2_s, lay6_fa2_c);
wire lay6_fa3_s, lay6_fa3_c;
full_adder lay6_fa3(lay6_fa2_s, lay5_ha0_c, lay5_fa3_c, lay6_fa3_s, lay6_fa3_c);
wire lay6_fa4_s, lay6_fa4_c;
full_adder lay6_fa4(lay6_fa3_s, lay5_fa2_c, lay5_fa1_c, lay6_fa4_s, lay6_fa4_c);
wire lay6_ha0_s, lay6_ha0_c;
half_adder lay6_ha0(lay6_fa4_s, lay5_fa0_c, lay6_ha0_s, lay6_ha0_c);
assign prod[6] = lay6_ha0_s;

wire lay7_fa0_s, lay7_fa0_c;
full_adder lay7_fa0(a7b0, a6b1, a5b2, lay7_fa0_s, lay7_fa0_c);
wire lay7_fa1_s, lay7_fa1_c;
full_adder lay7_fa1(lay7_fa0_s, a4b3, a3b4, lay7_fa1_s, lay7_fa1_c);
wire lay7_fa2_s, lay7_fa2_c;
full_adder lay7_fa2(lay7_fa1_s, a2b5, a1b6, lay7_fa2_s, lay7_fa2_c);
wire lay7_fa3_s, lay7_fa3_c;
full_adder lay7_fa3(lay7_fa2_s, a0b7, lay6_ha0_c, lay7_fa3_s, lay7_fa3_c);
wire lay7_fa4_s, lay7_fa4_c;
full_adder lay7_fa4(lay7_fa3_s, lay6_fa4_c, lay6_fa3_c, lay7_fa4_s, lay7_fa4_c);
wire lay7_fa5_s, lay7_fa5_c;
full_adder lay7_fa5(lay7_fa4_s, lay6_fa2_c, lay6_fa1_c, lay7_fa5_s, lay7_fa5_c);
wire lay7_ha0_s, lay7_ha0_c;
half_adder lay7_ha0(lay7_fa5_s, lay6_fa0_c, lay7_ha0_s, lay7_ha0_c);
assign prod[7] = lay7_ha0_s;

wire lay8_fa0_s, lay8_fa0_c;
full_adder lay8_fa0(a8b0, a7b1, a6b2, lay8_fa0_s, lay8_fa0_c);
wire lay8_fa1_s, lay8_fa1_c;
full_adder lay8_fa1(lay8_fa0_s, a5b3, a4b4, lay8_fa1_s, lay8_fa1_c);
wire lay8_fa2_s, lay8_fa2_c;
full_adder lay8_fa2(lay8_fa1_s, a3b5, a2b6, lay8_fa2_s, lay8_fa2_c);
wire lay8_fa3_s, lay8_fa3_c;
full_adder lay8_fa3(lay8_fa2_s, a1b7, a0b8, lay8_fa3_s, lay8_fa3_c);
wire lay8_fa4_s, lay8_fa4_c;
full_adder lay8_fa4(lay8_fa3_s, lay7_ha0_c, lay7_fa5_c, lay8_fa4_s, lay8_fa4_c);
wire lay8_fa5_s, lay8_fa5_c;
full_adder lay8_fa5(lay8_fa4_s, lay7_fa4_c, lay7_fa3_c, lay8_fa5_s, lay8_fa5_c);
wire lay8_fa6_s, lay8_fa6_c;
full_adder lay8_fa6(lay8_fa5_s, lay7_fa2_c, lay7_fa1_c, lay8_fa6_s, lay8_fa6_c);
wire lay8_ha0_s, lay8_ha0_c;
half_adder lay8_ha0(lay8_fa6_s, lay7_fa0_c, lay8_ha0_s, lay8_ha0_c);
assign prod[8] = lay8_ha0_s;

wire lay9_fa0_s, lay9_fa0_c;
full_adder lay9_fa0(a9b0, a8b1, a7b2, lay9_fa0_s, lay9_fa0_c);
wire lay9_fa1_s, lay9_fa1_c;
full_adder lay9_fa1(lay9_fa0_s, a6b3, a5b4, lay9_fa1_s, lay9_fa1_c);
wire lay9_fa2_s, lay9_fa2_c;
full_adder lay9_fa2(lay9_fa1_s, a4b5, a3b6, lay9_fa2_s, lay9_fa2_c);
wire lay9_fa3_s, lay9_fa3_c;
full_adder lay9_fa3(lay9_fa2_s, a2b7, a1b8, lay9_fa3_s, lay9_fa3_c);
wire lay9_fa4_s, lay9_fa4_c;
full_adder lay9_fa4(lay9_fa3_s, a0b9, lay8_ha0_c, lay9_fa4_s, lay9_fa4_c);
wire lay9_fa5_s, lay9_fa5_c;
full_adder lay9_fa5(lay9_fa4_s, lay8_fa6_c, lay8_fa5_c, lay9_fa5_s, lay9_fa5_c);
wire lay9_fa6_s, lay9_fa6_c;
full_adder lay9_fa6(lay9_fa5_s, lay8_fa4_c, lay8_fa3_c, lay9_fa6_s, lay9_fa6_c);
wire lay9_fa7_s, lay9_fa7_c;
full_adder lay9_fa7(lay9_fa6_s, lay8_fa2_c, lay8_fa1_c, lay9_fa7_s, lay9_fa7_c);
wire lay9_ha0_s, lay9_ha0_c;
half_adder lay9_ha0(lay9_fa7_s, lay8_fa0_c, lay9_ha0_s, lay9_ha0_c);
assign prod[9] = lay9_ha0_s;

wire lay10_fa0_s, lay10_fa0_c;
full_adder lay10_fa0(a10b0, a9b1, a8b2, lay10_fa0_s, lay10_fa0_c);
wire lay10_fa1_s, lay10_fa1_c;
full_adder lay10_fa1(lay10_fa0_s, a7b3, a6b4, lay10_fa1_s, lay10_fa1_c);
wire lay10_fa2_s, lay10_fa2_c;
full_adder lay10_fa2(lay10_fa1_s, a5b5, a4b6, lay10_fa2_s, lay10_fa2_c);
wire lay10_fa3_s, lay10_fa3_c;
full_adder lay10_fa3(lay10_fa2_s, a3b7, a2b8, lay10_fa3_s, lay10_fa3_c);
wire lay10_fa4_s, lay10_fa4_c;
full_adder lay10_fa4(lay10_fa3_s, a1b9, a0b10, lay10_fa4_s, lay10_fa4_c);
wire lay10_fa5_s, lay10_fa5_c;
full_adder lay10_fa5(lay10_fa4_s, lay9_ha0_c, lay9_fa7_c, lay10_fa5_s, lay10_fa5_c);
wire lay10_fa6_s, lay10_fa6_c;
full_adder lay10_fa6(lay10_fa5_s, lay9_fa6_c, lay9_fa5_c, lay10_fa6_s, lay10_fa6_c);
wire lay10_fa7_s, lay10_fa7_c;
full_adder lay10_fa7(lay10_fa6_s, lay9_fa4_c, lay9_fa3_c, lay10_fa7_s, lay10_fa7_c);
wire lay10_fa8_s, lay10_fa8_c;
full_adder lay10_fa8(lay10_fa7_s, lay9_fa2_c, lay9_fa1_c, lay10_fa8_s, lay10_fa8_c);
wire lay10_ha0_s, lay10_ha0_c;
half_adder lay10_ha0(lay10_fa8_s, lay9_fa0_c, lay10_ha0_s, lay10_ha0_c);
assign prod[10] = lay10_ha0_s;

wire lay11_fa0_s, lay11_fa0_c;
full_adder lay11_fa0(a11b0, a10b1, a9b2, lay11_fa0_s, lay11_fa0_c);
wire lay11_fa1_s, lay11_fa1_c;
full_adder lay11_fa1(lay11_fa0_s, a8b3, a7b4, lay11_fa1_s, lay11_fa1_c);
wire lay11_fa2_s, lay11_fa2_c;
full_adder lay11_fa2(lay11_fa1_s, a6b5, a5b6, lay11_fa2_s, lay11_fa2_c);
wire lay11_fa3_s, lay11_fa3_c;
full_adder lay11_fa3(lay11_fa2_s, a4b7, a3b8, lay11_fa3_s, lay11_fa3_c);
wire lay11_fa4_s, lay11_fa4_c;
full_adder lay11_fa4(lay11_fa3_s, a2b9, a1b10, lay11_fa4_s, lay11_fa4_c);
wire lay11_fa5_s, lay11_fa5_c;
full_adder lay11_fa5(lay11_fa4_s, a0b11, lay10_ha0_c, lay11_fa5_s, lay11_fa5_c);
wire lay11_fa6_s, lay11_fa6_c;
full_adder lay11_fa6(lay11_fa5_s, lay10_fa8_c, lay10_fa7_c, lay11_fa6_s, lay11_fa6_c);
wire lay11_fa7_s, lay11_fa7_c;
full_adder lay11_fa7(lay11_fa6_s, lay10_fa6_c, lay10_fa5_c, lay11_fa7_s, lay11_fa7_c);
wire lay11_fa8_s, lay11_fa8_c;
full_adder lay11_fa8(lay11_fa7_s, lay10_fa4_c, lay10_fa3_c, lay11_fa8_s, lay11_fa8_c);
wire lay11_fa9_s, lay11_fa9_c;
full_adder lay11_fa9(lay11_fa8_s, lay10_fa2_c, lay10_fa1_c, lay11_fa9_s, lay11_fa9_c);
wire lay11_ha0_s, lay11_ha0_c;
half_adder lay11_ha0(lay11_fa9_s, lay10_fa0_c, lay11_ha0_s, lay11_ha0_c);
assign prod[11] = lay11_ha0_s;

wire lay12_fa0_s, lay12_fa0_c;
full_adder lay12_fa0(a12b0, a11b1, a10b2, lay12_fa0_s, lay12_fa0_c);
wire lay12_fa1_s, lay12_fa1_c;
full_adder lay12_fa1(lay12_fa0_s, a9b3, a8b4, lay12_fa1_s, lay12_fa1_c);
wire lay12_fa2_s, lay12_fa2_c;
full_adder lay12_fa2(lay12_fa1_s, a7b5, a6b6, lay12_fa2_s, lay12_fa2_c);
wire lay12_fa3_s, lay12_fa3_c;
full_adder lay12_fa3(lay12_fa2_s, a5b7, a4b8, lay12_fa3_s, lay12_fa3_c);
wire lay12_fa4_s, lay12_fa4_c;
full_adder lay12_fa4(lay12_fa3_s, a3b9, a2b10, lay12_fa4_s, lay12_fa4_c);
wire lay12_fa5_s, lay12_fa5_c;
full_adder lay12_fa5(lay12_fa4_s, a1b11, a0b12, lay12_fa5_s, lay12_fa5_c);
wire lay12_fa6_s, lay12_fa6_c;
full_adder lay12_fa6(lay12_fa5_s, lay11_ha0_c, lay11_fa9_c, lay12_fa6_s, lay12_fa6_c);
wire lay12_fa7_s, lay12_fa7_c;
full_adder lay12_fa7(lay12_fa6_s, lay11_fa8_c, lay11_fa7_c, lay12_fa7_s, lay12_fa7_c);
wire lay12_fa8_s, lay12_fa8_c;
full_adder lay12_fa8(lay12_fa7_s, lay11_fa6_c, lay11_fa5_c, lay12_fa8_s, lay12_fa8_c);
wire lay12_fa9_s, lay12_fa9_c;
full_adder lay12_fa9(lay12_fa8_s, lay11_fa4_c, lay11_fa3_c, lay12_fa9_s, lay12_fa9_c);
wire lay12_fa10_s, lay12_fa10_c;
full_adder lay12_fa10(lay12_fa9_s, lay11_fa2_c, lay11_fa1_c, lay12_fa10_s, lay12_fa10_c);
wire lay12_ha0_s, lay12_ha0_c;
half_adder lay12_ha0(lay12_fa10_s, lay11_fa0_c, lay12_ha0_s, lay12_ha0_c);
assign prod[12] = lay12_ha0_s;

wire lay13_fa0_s, lay13_fa0_c;
full_adder lay13_fa0(a13b0, a12b1, a11b2, lay13_fa0_s, lay13_fa0_c);
wire lay13_fa1_s, lay13_fa1_c;
full_adder lay13_fa1(lay13_fa0_s, a10b3, a9b4, lay13_fa1_s, lay13_fa1_c);
wire lay13_fa2_s, lay13_fa2_c;
full_adder lay13_fa2(lay13_fa1_s, a8b5, a7b6, lay13_fa2_s, lay13_fa2_c);
wire lay13_fa3_s, lay13_fa3_c;
full_adder lay13_fa3(lay13_fa2_s, a6b7, a5b8, lay13_fa3_s, lay13_fa3_c);
wire lay13_fa4_s, lay13_fa4_c;
full_adder lay13_fa4(lay13_fa3_s, a4b9, a3b10, lay13_fa4_s, lay13_fa4_c);
wire lay13_fa5_s, lay13_fa5_c;
full_adder lay13_fa5(lay13_fa4_s, a2b11, a1b12, lay13_fa5_s, lay13_fa5_c);
wire lay13_fa6_s, lay13_fa6_c;
full_adder lay13_fa6(lay13_fa5_s, a0b13, lay12_ha0_c, lay13_fa6_s, lay13_fa6_c);
wire lay13_fa7_s, lay13_fa7_c;
full_adder lay13_fa7(lay13_fa6_s, lay12_fa10_c, lay12_fa9_c, lay13_fa7_s, lay13_fa7_c);
wire lay13_fa8_s, lay13_fa8_c;
full_adder lay13_fa8(lay13_fa7_s, lay12_fa8_c, lay12_fa7_c, lay13_fa8_s, lay13_fa8_c);
wire lay13_fa9_s, lay13_fa9_c;
full_adder lay13_fa9(lay13_fa8_s, lay12_fa6_c, lay12_fa5_c, lay13_fa9_s, lay13_fa9_c);
wire lay13_fa10_s, lay13_fa10_c;
full_adder lay13_fa10(lay13_fa9_s, lay12_fa4_c, lay12_fa3_c, lay13_fa10_s, lay13_fa10_c);
wire lay13_fa11_s, lay13_fa11_c;
full_adder lay13_fa11(lay13_fa10_s, lay12_fa2_c, lay12_fa1_c, lay13_fa11_s, lay13_fa11_c);
wire lay13_ha0_s, lay13_ha0_c;
half_adder lay13_ha0(lay13_fa11_s, lay12_fa0_c, lay13_ha0_s, lay13_ha0_c);
assign prod[13] = lay13_ha0_s;

wire lay14_fa0_s, lay14_fa0_c;
full_adder lay14_fa0(a14b0, a13b1, a12b2, lay14_fa0_s, lay14_fa0_c);
wire lay14_fa1_s, lay14_fa1_c;
full_adder lay14_fa1(lay14_fa0_s, a11b3, a10b4, lay14_fa1_s, lay14_fa1_c);
wire lay14_fa2_s, lay14_fa2_c;
full_adder lay14_fa2(lay14_fa1_s, a9b5, a8b6, lay14_fa2_s, lay14_fa2_c);
wire lay14_fa3_s, lay14_fa3_c;
full_adder lay14_fa3(lay14_fa2_s, a7b7, a6b8, lay14_fa3_s, lay14_fa3_c);
wire lay14_fa4_s, lay14_fa4_c;
full_adder lay14_fa4(lay14_fa3_s, a5b9, a4b10, lay14_fa4_s, lay14_fa4_c);
wire lay14_fa5_s, lay14_fa5_c;
full_adder lay14_fa5(lay14_fa4_s, a3b11, a2b12, lay14_fa5_s, lay14_fa5_c);
wire lay14_fa6_s, lay14_fa6_c;
full_adder lay14_fa6(lay14_fa5_s, a1b13, a0b14, lay14_fa6_s, lay14_fa6_c);
wire lay14_fa7_s, lay14_fa7_c;
full_adder lay14_fa7(lay14_fa6_s, lay13_ha0_c, lay13_fa11_c, lay14_fa7_s, lay14_fa7_c);
wire lay14_fa8_s, lay14_fa8_c;
full_adder lay14_fa8(lay14_fa7_s, lay13_fa10_c, lay13_fa9_c, lay14_fa8_s, lay14_fa8_c);
wire lay14_fa9_s, lay14_fa9_c;
full_adder lay14_fa9(lay14_fa8_s, lay13_fa8_c, lay13_fa7_c, lay14_fa9_s, lay14_fa9_c);
wire lay14_fa10_s, lay14_fa10_c;
full_adder lay14_fa10(lay14_fa9_s, lay13_fa6_c, lay13_fa5_c, lay14_fa10_s, lay14_fa10_c);
wire lay14_fa11_s, lay14_fa11_c;
full_adder lay14_fa11(lay14_fa10_s, lay13_fa4_c, lay13_fa3_c, lay14_fa11_s, lay14_fa11_c);
wire lay14_fa12_s, lay14_fa12_c;
full_adder lay14_fa12(lay14_fa11_s, lay13_fa2_c, lay13_fa1_c, lay14_fa12_s, lay14_fa12_c);
wire lay14_ha0_s, lay14_ha0_c;
half_adder lay14_ha0(lay14_fa12_s, lay13_fa0_c, lay14_ha0_s, lay14_ha0_c);
assign prod[14] = lay14_ha0_s;

wire lay15_fa0_s, lay15_fa0_c;
full_adder lay15_fa0(a15b0, a14b1, a13b2, lay15_fa0_s, lay15_fa0_c);
wire lay15_fa1_s, lay15_fa1_c;
full_adder lay15_fa1(lay15_fa0_s, a12b3, a11b4, lay15_fa1_s, lay15_fa1_c);
wire lay15_fa2_s, lay15_fa2_c;
full_adder lay15_fa2(lay15_fa1_s, a10b5, a9b6, lay15_fa2_s, lay15_fa2_c);
wire lay15_fa3_s, lay15_fa3_c;
full_adder lay15_fa3(lay15_fa2_s, a8b7, a7b8, lay15_fa3_s, lay15_fa3_c);
wire lay15_fa4_s, lay15_fa4_c;
full_adder lay15_fa4(lay15_fa3_s, a6b9, a5b10, lay15_fa4_s, lay15_fa4_c);
wire lay15_fa5_s, lay15_fa5_c;
full_adder lay15_fa5(lay15_fa4_s, a4b11, a3b12, lay15_fa5_s, lay15_fa5_c);
wire lay15_fa6_s, lay15_fa6_c;
full_adder lay15_fa6(lay15_fa5_s, a2b13, a1b14, lay15_fa6_s, lay15_fa6_c);
wire lay15_fa7_s, lay15_fa7_c;
full_adder lay15_fa7(lay15_fa6_s, a0b15, lay14_ha0_c, lay15_fa7_s, lay15_fa7_c);
wire lay15_fa8_s, lay15_fa8_c;
full_adder lay15_fa8(lay15_fa7_s, lay14_fa12_c, lay14_fa11_c, lay15_fa8_s, lay15_fa8_c);
wire lay15_fa9_s, lay15_fa9_c;
full_adder lay15_fa9(lay15_fa8_s, lay14_fa10_c, lay14_fa9_c, lay15_fa9_s, lay15_fa9_c);
wire lay15_fa10_s, lay15_fa10_c;
full_adder lay15_fa10(lay15_fa9_s, lay14_fa8_c, lay14_fa7_c, lay15_fa10_s, lay15_fa10_c);
wire lay15_fa11_s, lay15_fa11_c;
full_adder lay15_fa11(lay15_fa10_s, lay14_fa6_c, lay14_fa5_c, lay15_fa11_s, lay15_fa11_c);
wire lay15_fa12_s, lay15_fa12_c;
full_adder lay15_fa12(lay15_fa11_s, lay14_fa4_c, lay14_fa3_c, lay15_fa12_s, lay15_fa12_c);
wire lay15_fa13_s, lay15_fa13_c;
full_adder lay15_fa13(lay15_fa12_s, lay14_fa2_c, lay14_fa1_c, lay15_fa13_s, lay15_fa13_c);
wire lay15_ha0_s, lay15_ha0_c;
half_adder lay15_ha0(lay15_fa13_s, lay14_fa0_c, lay15_ha0_s, lay15_ha0_c);
assign prod[15] = lay15_ha0_s;

wire lay16_fa0_s, lay16_fa0_c;
full_adder lay16_fa0(a16b0, a15b1, a14b2, lay16_fa0_s, lay16_fa0_c);
wire lay16_fa1_s, lay16_fa1_c;
full_adder lay16_fa1(lay16_fa0_s, a13b3, a12b4, lay16_fa1_s, lay16_fa1_c);
wire lay16_fa2_s, lay16_fa2_c;
full_adder lay16_fa2(lay16_fa1_s, a11b5, a10b6, lay16_fa2_s, lay16_fa2_c);
wire lay16_fa3_s, lay16_fa3_c;
full_adder lay16_fa3(lay16_fa2_s, a9b7, a8b8, lay16_fa3_s, lay16_fa3_c);
wire lay16_fa4_s, lay16_fa4_c;
full_adder lay16_fa4(lay16_fa3_s, a7b9, a6b10, lay16_fa4_s, lay16_fa4_c);
wire lay16_fa5_s, lay16_fa5_c;
full_adder lay16_fa5(lay16_fa4_s, a5b11, a4b12, lay16_fa5_s, lay16_fa5_c);
wire lay16_fa6_s, lay16_fa6_c;
full_adder lay16_fa6(lay16_fa5_s, a3b13, a2b14, lay16_fa6_s, lay16_fa6_c);
wire lay16_fa7_s, lay16_fa7_c;
full_adder lay16_fa7(lay16_fa6_s, a1b15, a0b16, lay16_fa7_s, lay16_fa7_c);
wire lay16_fa8_s, lay16_fa8_c;
full_adder lay16_fa8(lay16_fa7_s, lay15_ha0_c, lay15_fa13_c, lay16_fa8_s, lay16_fa8_c);
wire lay16_fa9_s, lay16_fa9_c;
full_adder lay16_fa9(lay16_fa8_s, lay15_fa12_c, lay15_fa11_c, lay16_fa9_s, lay16_fa9_c);
wire lay16_fa10_s, lay16_fa10_c;
full_adder lay16_fa10(lay16_fa9_s, lay15_fa10_c, lay15_fa9_c, lay16_fa10_s, lay16_fa10_c);
wire lay16_fa11_s, lay16_fa11_c;
full_adder lay16_fa11(lay16_fa10_s, lay15_fa8_c, lay15_fa7_c, lay16_fa11_s, lay16_fa11_c);
wire lay16_fa12_s, lay16_fa12_c;
full_adder lay16_fa12(lay16_fa11_s, lay15_fa6_c, lay15_fa5_c, lay16_fa12_s, lay16_fa12_c);
wire lay16_fa13_s, lay16_fa13_c;
full_adder lay16_fa13(lay16_fa12_s, lay15_fa4_c, lay15_fa3_c, lay16_fa13_s, lay16_fa13_c);
wire lay16_fa14_s, lay16_fa14_c;
full_adder lay16_fa14(lay16_fa13_s, lay15_fa2_c, lay15_fa1_c, lay16_fa14_s, lay16_fa14_c);
wire lay16_ha0_s, lay16_ha0_c;
half_adder lay16_ha0(lay16_fa14_s, lay15_fa0_c, lay16_ha0_s, lay16_ha0_c);
assign prod[16] = lay16_ha0_s;

wire lay17_fa0_s, lay17_fa0_c;
full_adder lay17_fa0(a17b0, a16b1, a15b2, lay17_fa0_s, lay17_fa0_c);
wire lay17_fa1_s, lay17_fa1_c;
full_adder lay17_fa1(lay17_fa0_s, a14b3, a13b4, lay17_fa1_s, lay17_fa1_c);
wire lay17_fa2_s, lay17_fa2_c;
full_adder lay17_fa2(lay17_fa1_s, a12b5, a11b6, lay17_fa2_s, lay17_fa2_c);
wire lay17_fa3_s, lay17_fa3_c;
full_adder lay17_fa3(lay17_fa2_s, a10b7, a9b8, lay17_fa3_s, lay17_fa3_c);
wire lay17_fa4_s, lay17_fa4_c;
full_adder lay17_fa4(lay17_fa3_s, a8b9, a7b10, lay17_fa4_s, lay17_fa4_c);
wire lay17_fa5_s, lay17_fa5_c;
full_adder lay17_fa5(lay17_fa4_s, a6b11, a5b12, lay17_fa5_s, lay17_fa5_c);
wire lay17_fa6_s, lay17_fa6_c;
full_adder lay17_fa6(lay17_fa5_s, a4b13, a3b14, lay17_fa6_s, lay17_fa6_c);
wire lay17_fa7_s, lay17_fa7_c;
full_adder lay17_fa7(lay17_fa6_s, a2b15, a1b16, lay17_fa7_s, lay17_fa7_c);
wire lay17_fa8_s, lay17_fa8_c;
full_adder lay17_fa8(lay17_fa7_s, a0b17, lay16_ha0_c, lay17_fa8_s, lay17_fa8_c);
wire lay17_fa9_s, lay17_fa9_c;
full_adder lay17_fa9(lay17_fa8_s, lay16_fa14_c, lay16_fa13_c, lay17_fa9_s, lay17_fa9_c);
wire lay17_fa10_s, lay17_fa10_c;
full_adder lay17_fa10(lay17_fa9_s, lay16_fa12_c, lay16_fa11_c, lay17_fa10_s, lay17_fa10_c);
wire lay17_fa11_s, lay17_fa11_c;
full_adder lay17_fa11(lay17_fa10_s, lay16_fa10_c, lay16_fa9_c, lay17_fa11_s, lay17_fa11_c);
wire lay17_fa12_s, lay17_fa12_c;
full_adder lay17_fa12(lay17_fa11_s, lay16_fa8_c, lay16_fa7_c, lay17_fa12_s, lay17_fa12_c);
wire lay17_fa13_s, lay17_fa13_c;
full_adder lay17_fa13(lay17_fa12_s, lay16_fa6_c, lay16_fa5_c, lay17_fa13_s, lay17_fa13_c);
wire lay17_fa14_s, lay17_fa14_c;
full_adder lay17_fa14(lay17_fa13_s, lay16_fa4_c, lay16_fa3_c, lay17_fa14_s, lay17_fa14_c);
wire lay17_fa15_s, lay17_fa15_c;
full_adder lay17_fa15(lay17_fa14_s, lay16_fa2_c, lay16_fa1_c, lay17_fa15_s, lay17_fa15_c);
wire lay17_ha0_s, lay17_ha0_c;
half_adder lay17_ha0(lay17_fa15_s, lay16_fa0_c, lay17_ha0_s, lay17_ha0_c);
assign prod[17] = lay17_ha0_s;

wire lay18_fa0_s, lay18_fa0_c;
full_adder lay18_fa0(a18b0, a17b1, a16b2, lay18_fa0_s, lay18_fa0_c);
wire lay18_fa1_s, lay18_fa1_c;
full_adder lay18_fa1(lay18_fa0_s, a15b3, a14b4, lay18_fa1_s, lay18_fa1_c);
wire lay18_fa2_s, lay18_fa2_c;
full_adder lay18_fa2(lay18_fa1_s, a13b5, a12b6, lay18_fa2_s, lay18_fa2_c);
wire lay18_fa3_s, lay18_fa3_c;
full_adder lay18_fa3(lay18_fa2_s, a11b7, a10b8, lay18_fa3_s, lay18_fa3_c);
wire lay18_fa4_s, lay18_fa4_c;
full_adder lay18_fa4(lay18_fa3_s, a9b9, a8b10, lay18_fa4_s, lay18_fa4_c);
wire lay18_fa5_s, lay18_fa5_c;
full_adder lay18_fa5(lay18_fa4_s, a7b11, a6b12, lay18_fa5_s, lay18_fa5_c);
wire lay18_fa6_s, lay18_fa6_c;
full_adder lay18_fa6(lay18_fa5_s, a5b13, a4b14, lay18_fa6_s, lay18_fa6_c);
wire lay18_fa7_s, lay18_fa7_c;
full_adder lay18_fa7(lay18_fa6_s, a3b15, a2b16, lay18_fa7_s, lay18_fa7_c);
wire lay18_fa8_s, lay18_fa8_c;
full_adder lay18_fa8(lay18_fa7_s, a1b17, a0b18, lay18_fa8_s, lay18_fa8_c);
wire lay18_fa9_s, lay18_fa9_c;
full_adder lay18_fa9(lay18_fa8_s, lay17_ha0_c, lay17_fa15_c, lay18_fa9_s, lay18_fa9_c);
wire lay18_fa10_s, lay18_fa10_c;
full_adder lay18_fa10(lay18_fa9_s, lay17_fa14_c, lay17_fa13_c, lay18_fa10_s, lay18_fa10_c);
wire lay18_fa11_s, lay18_fa11_c;
full_adder lay18_fa11(lay18_fa10_s, lay17_fa12_c, lay17_fa11_c, lay18_fa11_s, lay18_fa11_c);
wire lay18_fa12_s, lay18_fa12_c;
full_adder lay18_fa12(lay18_fa11_s, lay17_fa10_c, lay17_fa9_c, lay18_fa12_s, lay18_fa12_c);
wire lay18_fa13_s, lay18_fa13_c;
full_adder lay18_fa13(lay18_fa12_s, lay17_fa8_c, lay17_fa7_c, lay18_fa13_s, lay18_fa13_c);
wire lay18_fa14_s, lay18_fa14_c;
full_adder lay18_fa14(lay18_fa13_s, lay17_fa6_c, lay17_fa5_c, lay18_fa14_s, lay18_fa14_c);
wire lay18_fa15_s, lay18_fa15_c;
full_adder lay18_fa15(lay18_fa14_s, lay17_fa4_c, lay17_fa3_c, lay18_fa15_s, lay18_fa15_c);
wire lay18_fa16_s, lay18_fa16_c;
full_adder lay18_fa16(lay18_fa15_s, lay17_fa2_c, lay17_fa1_c, lay18_fa16_s, lay18_fa16_c);
wire lay18_ha0_s, lay18_ha0_c;
half_adder lay18_ha0(lay18_fa16_s, lay17_fa0_c, lay18_ha0_s, lay18_ha0_c);
assign prod[18] = lay18_ha0_s;

wire lay19_fa0_s, lay19_fa0_c;
full_adder lay19_fa0(a19b0, a18b1, a17b2, lay19_fa0_s, lay19_fa0_c);
wire lay19_fa1_s, lay19_fa1_c;
full_adder lay19_fa1(lay19_fa0_s, a16b3, a15b4, lay19_fa1_s, lay19_fa1_c);
wire lay19_fa2_s, lay19_fa2_c;
full_adder lay19_fa2(lay19_fa1_s, a14b5, a13b6, lay19_fa2_s, lay19_fa2_c);
wire lay19_fa3_s, lay19_fa3_c;
full_adder lay19_fa3(lay19_fa2_s, a12b7, a11b8, lay19_fa3_s, lay19_fa3_c);
wire lay19_fa4_s, lay19_fa4_c;
full_adder lay19_fa4(lay19_fa3_s, a10b9, a9b10, lay19_fa4_s, lay19_fa4_c);
wire lay19_fa5_s, lay19_fa5_c;
full_adder lay19_fa5(lay19_fa4_s, a8b11, a7b12, lay19_fa5_s, lay19_fa5_c);
wire lay19_fa6_s, lay19_fa6_c;
full_adder lay19_fa6(lay19_fa5_s, a6b13, a5b14, lay19_fa6_s, lay19_fa6_c);
wire lay19_fa7_s, lay19_fa7_c;
full_adder lay19_fa7(lay19_fa6_s, a4b15, a3b16, lay19_fa7_s, lay19_fa7_c);
wire lay19_fa8_s, lay19_fa8_c;
full_adder lay19_fa8(lay19_fa7_s, a2b17, a1b18, lay19_fa8_s, lay19_fa8_c);
wire lay19_fa9_s, lay19_fa9_c;
full_adder lay19_fa9(lay19_fa8_s, a0b19, lay18_ha0_c, lay19_fa9_s, lay19_fa9_c);
wire lay19_fa10_s, lay19_fa10_c;
full_adder lay19_fa10(lay19_fa9_s, lay18_fa16_c, lay18_fa15_c, lay19_fa10_s, lay19_fa10_c);
wire lay19_fa11_s, lay19_fa11_c;
full_adder lay19_fa11(lay19_fa10_s, lay18_fa14_c, lay18_fa13_c, lay19_fa11_s, lay19_fa11_c);
wire lay19_fa12_s, lay19_fa12_c;
full_adder lay19_fa12(lay19_fa11_s, lay18_fa12_c, lay18_fa11_c, lay19_fa12_s, lay19_fa12_c);
wire lay19_fa13_s, lay19_fa13_c;
full_adder lay19_fa13(lay19_fa12_s, lay18_fa10_c, lay18_fa9_c, lay19_fa13_s, lay19_fa13_c);
wire lay19_fa14_s, lay19_fa14_c;
full_adder lay19_fa14(lay19_fa13_s, lay18_fa8_c, lay18_fa7_c, lay19_fa14_s, lay19_fa14_c);
wire lay19_fa15_s, lay19_fa15_c;
full_adder lay19_fa15(lay19_fa14_s, lay18_fa6_c, lay18_fa5_c, lay19_fa15_s, lay19_fa15_c);
wire lay19_fa16_s, lay19_fa16_c;
full_adder lay19_fa16(lay19_fa15_s, lay18_fa4_c, lay18_fa3_c, lay19_fa16_s, lay19_fa16_c);
wire lay19_fa17_s, lay19_fa17_c;
full_adder lay19_fa17(lay19_fa16_s, lay18_fa2_c, lay18_fa1_c, lay19_fa17_s, lay19_fa17_c);
wire lay19_ha0_s, lay19_ha0_c;
half_adder lay19_ha0(lay19_fa17_s, lay18_fa0_c, lay19_ha0_s, lay19_ha0_c);
assign prod[19] = lay19_ha0_s;

wire lay20_fa0_s, lay20_fa0_c;
full_adder lay20_fa0(a20b0, a19b1, a18b2, lay20_fa0_s, lay20_fa0_c);
wire lay20_fa1_s, lay20_fa1_c;
full_adder lay20_fa1(lay20_fa0_s, a17b3, a16b4, lay20_fa1_s, lay20_fa1_c);
wire lay20_fa2_s, lay20_fa2_c;
full_adder lay20_fa2(lay20_fa1_s, a15b5, a14b6, lay20_fa2_s, lay20_fa2_c);
wire lay20_fa3_s, lay20_fa3_c;
full_adder lay20_fa3(lay20_fa2_s, a13b7, a12b8, lay20_fa3_s, lay20_fa3_c);
wire lay20_fa4_s, lay20_fa4_c;
full_adder lay20_fa4(lay20_fa3_s, a11b9, a10b10, lay20_fa4_s, lay20_fa4_c);
wire lay20_fa5_s, lay20_fa5_c;
full_adder lay20_fa5(lay20_fa4_s, a9b11, a8b12, lay20_fa5_s, lay20_fa5_c);
wire lay20_fa6_s, lay20_fa6_c;
full_adder lay20_fa6(lay20_fa5_s, a7b13, a6b14, lay20_fa6_s, lay20_fa6_c);
wire lay20_fa7_s, lay20_fa7_c;
full_adder lay20_fa7(lay20_fa6_s, a5b15, a4b16, lay20_fa7_s, lay20_fa7_c);
wire lay20_fa8_s, lay20_fa8_c;
full_adder lay20_fa8(lay20_fa7_s, a3b17, a2b18, lay20_fa8_s, lay20_fa8_c);
wire lay20_fa9_s, lay20_fa9_c;
full_adder lay20_fa9(lay20_fa8_s, a1b19, a0b20, lay20_fa9_s, lay20_fa9_c);
wire lay20_fa10_s, lay20_fa10_c;
full_adder lay20_fa10(lay20_fa9_s, lay19_ha0_c, lay19_fa17_c, lay20_fa10_s, lay20_fa10_c);
wire lay20_fa11_s, lay20_fa11_c;
full_adder lay20_fa11(lay20_fa10_s, lay19_fa16_c, lay19_fa15_c, lay20_fa11_s, lay20_fa11_c);
wire lay20_fa12_s, lay20_fa12_c;
full_adder lay20_fa12(lay20_fa11_s, lay19_fa14_c, lay19_fa13_c, lay20_fa12_s, lay20_fa12_c);
wire lay20_fa13_s, lay20_fa13_c;
full_adder lay20_fa13(lay20_fa12_s, lay19_fa12_c, lay19_fa11_c, lay20_fa13_s, lay20_fa13_c);
wire lay20_fa14_s, lay20_fa14_c;
full_adder lay20_fa14(lay20_fa13_s, lay19_fa10_c, lay19_fa9_c, lay20_fa14_s, lay20_fa14_c);
wire lay20_fa15_s, lay20_fa15_c;
full_adder lay20_fa15(lay20_fa14_s, lay19_fa8_c, lay19_fa7_c, lay20_fa15_s, lay20_fa15_c);
wire lay20_fa16_s, lay20_fa16_c;
full_adder lay20_fa16(lay20_fa15_s, lay19_fa6_c, lay19_fa5_c, lay20_fa16_s, lay20_fa16_c);
wire lay20_fa17_s, lay20_fa17_c;
full_adder lay20_fa17(lay20_fa16_s, lay19_fa4_c, lay19_fa3_c, lay20_fa17_s, lay20_fa17_c);
wire lay20_fa18_s, lay20_fa18_c;
full_adder lay20_fa18(lay20_fa17_s, lay19_fa2_c, lay19_fa1_c, lay20_fa18_s, lay20_fa18_c);
wire lay20_ha0_s, lay20_ha0_c;
half_adder lay20_ha0(lay20_fa18_s, lay19_fa0_c, lay20_ha0_s, lay20_ha0_c);
assign prod[20] = lay20_ha0_s;

wire lay21_fa0_s, lay21_fa0_c;
full_adder lay21_fa0(a21b0, a20b1, a19b2, lay21_fa0_s, lay21_fa0_c);
wire lay21_fa1_s, lay21_fa1_c;
full_adder lay21_fa1(lay21_fa0_s, a18b3, a17b4, lay21_fa1_s, lay21_fa1_c);
wire lay21_fa2_s, lay21_fa2_c;
full_adder lay21_fa2(lay21_fa1_s, a16b5, a15b6, lay21_fa2_s, lay21_fa2_c);
wire lay21_fa3_s, lay21_fa3_c;
full_adder lay21_fa3(lay21_fa2_s, a14b7, a13b8, lay21_fa3_s, lay21_fa3_c);
wire lay21_fa4_s, lay21_fa4_c;
full_adder lay21_fa4(lay21_fa3_s, a12b9, a11b10, lay21_fa4_s, lay21_fa4_c);
wire lay21_fa5_s, lay21_fa5_c;
full_adder lay21_fa5(lay21_fa4_s, a10b11, a9b12, lay21_fa5_s, lay21_fa5_c);
wire lay21_fa6_s, lay21_fa6_c;
full_adder lay21_fa6(lay21_fa5_s, a8b13, a7b14, lay21_fa6_s, lay21_fa6_c);
wire lay21_fa7_s, lay21_fa7_c;
full_adder lay21_fa7(lay21_fa6_s, a6b15, a5b16, lay21_fa7_s, lay21_fa7_c);
wire lay21_fa8_s, lay21_fa8_c;
full_adder lay21_fa8(lay21_fa7_s, a4b17, a3b18, lay21_fa8_s, lay21_fa8_c);
wire lay21_fa9_s, lay21_fa9_c;
full_adder lay21_fa9(lay21_fa8_s, a2b19, a1b20, lay21_fa9_s, lay21_fa9_c);
wire lay21_fa10_s, lay21_fa10_c;
full_adder lay21_fa10(lay21_fa9_s, a0b21, lay20_ha0_c, lay21_fa10_s, lay21_fa10_c);
wire lay21_fa11_s, lay21_fa11_c;
full_adder lay21_fa11(lay21_fa10_s, lay20_fa18_c, lay20_fa17_c, lay21_fa11_s, lay21_fa11_c);
wire lay21_fa12_s, lay21_fa12_c;
full_adder lay21_fa12(lay21_fa11_s, lay20_fa16_c, lay20_fa15_c, lay21_fa12_s, lay21_fa12_c);
wire lay21_fa13_s, lay21_fa13_c;
full_adder lay21_fa13(lay21_fa12_s, lay20_fa14_c, lay20_fa13_c, lay21_fa13_s, lay21_fa13_c);
wire lay21_fa14_s, lay21_fa14_c;
full_adder lay21_fa14(lay21_fa13_s, lay20_fa12_c, lay20_fa11_c, lay21_fa14_s, lay21_fa14_c);
wire lay21_fa15_s, lay21_fa15_c;
full_adder lay21_fa15(lay21_fa14_s, lay20_fa10_c, lay20_fa9_c, lay21_fa15_s, lay21_fa15_c);
wire lay21_fa16_s, lay21_fa16_c;
full_adder lay21_fa16(lay21_fa15_s, lay20_fa8_c, lay20_fa7_c, lay21_fa16_s, lay21_fa16_c);
wire lay21_fa17_s, lay21_fa17_c;
full_adder lay21_fa17(lay21_fa16_s, lay20_fa6_c, lay20_fa5_c, lay21_fa17_s, lay21_fa17_c);
wire lay21_fa18_s, lay21_fa18_c;
full_adder lay21_fa18(lay21_fa17_s, lay20_fa4_c, lay20_fa3_c, lay21_fa18_s, lay21_fa18_c);
wire lay21_fa19_s, lay21_fa19_c;
full_adder lay21_fa19(lay21_fa18_s, lay20_fa2_c, lay20_fa1_c, lay21_fa19_s, lay21_fa19_c);
wire lay21_ha0_s, lay21_ha0_c;
half_adder lay21_ha0(lay21_fa19_s, lay20_fa0_c, lay21_ha0_s, lay21_ha0_c);
assign prod[21] = lay21_ha0_s;

wire lay22_fa0_s, lay22_fa0_c;
full_adder lay22_fa0(a22b0, a21b1, a20b2, lay22_fa0_s, lay22_fa0_c);
wire lay22_fa1_s, lay22_fa1_c;
full_adder lay22_fa1(lay22_fa0_s, a19b3, a18b4, lay22_fa1_s, lay22_fa1_c);
wire lay22_fa2_s, lay22_fa2_c;
full_adder lay22_fa2(lay22_fa1_s, a17b5, a16b6, lay22_fa2_s, lay22_fa2_c);
wire lay22_fa3_s, lay22_fa3_c;
full_adder lay22_fa3(lay22_fa2_s, a15b7, a14b8, lay22_fa3_s, lay22_fa3_c);
wire lay22_fa4_s, lay22_fa4_c;
full_adder lay22_fa4(lay22_fa3_s, a13b9, a12b10, lay22_fa4_s, lay22_fa4_c);
wire lay22_fa5_s, lay22_fa5_c;
full_adder lay22_fa5(lay22_fa4_s, a11b11, a10b12, lay22_fa5_s, lay22_fa5_c);
wire lay22_fa6_s, lay22_fa6_c;
full_adder lay22_fa6(lay22_fa5_s, a9b13, a8b14, lay22_fa6_s, lay22_fa6_c);
wire lay22_fa7_s, lay22_fa7_c;
full_adder lay22_fa7(lay22_fa6_s, a7b15, a6b16, lay22_fa7_s, lay22_fa7_c);
wire lay22_fa8_s, lay22_fa8_c;
full_adder lay22_fa8(lay22_fa7_s, a5b17, a4b18, lay22_fa8_s, lay22_fa8_c);
wire lay22_fa9_s, lay22_fa9_c;
full_adder lay22_fa9(lay22_fa8_s, a3b19, a2b20, lay22_fa9_s, lay22_fa9_c);
wire lay22_fa10_s, lay22_fa10_c;
full_adder lay22_fa10(lay22_fa9_s, a1b21, a0b22, lay22_fa10_s, lay22_fa10_c);
wire lay22_fa11_s, lay22_fa11_c;
full_adder lay22_fa11(lay22_fa10_s, lay21_ha0_c, lay21_fa19_c, lay22_fa11_s, lay22_fa11_c);
wire lay22_fa12_s, lay22_fa12_c;
full_adder lay22_fa12(lay22_fa11_s, lay21_fa18_c, lay21_fa17_c, lay22_fa12_s, lay22_fa12_c);
wire lay22_fa13_s, lay22_fa13_c;
full_adder lay22_fa13(lay22_fa12_s, lay21_fa16_c, lay21_fa15_c, lay22_fa13_s, lay22_fa13_c);
wire lay22_fa14_s, lay22_fa14_c;
full_adder lay22_fa14(lay22_fa13_s, lay21_fa14_c, lay21_fa13_c, lay22_fa14_s, lay22_fa14_c);
wire lay22_fa15_s, lay22_fa15_c;
full_adder lay22_fa15(lay22_fa14_s, lay21_fa12_c, lay21_fa11_c, lay22_fa15_s, lay22_fa15_c);
wire lay22_fa16_s, lay22_fa16_c;
full_adder lay22_fa16(lay22_fa15_s, lay21_fa10_c, lay21_fa9_c, lay22_fa16_s, lay22_fa16_c);
wire lay22_fa17_s, lay22_fa17_c;
full_adder lay22_fa17(lay22_fa16_s, lay21_fa8_c, lay21_fa7_c, lay22_fa17_s, lay22_fa17_c);
wire lay22_fa18_s, lay22_fa18_c;
full_adder lay22_fa18(lay22_fa17_s, lay21_fa6_c, lay21_fa5_c, lay22_fa18_s, lay22_fa18_c);
wire lay22_fa19_s, lay22_fa19_c;
full_adder lay22_fa19(lay22_fa18_s, lay21_fa4_c, lay21_fa3_c, lay22_fa19_s, lay22_fa19_c);
wire lay22_fa20_s, lay22_fa20_c;
full_adder lay22_fa20(lay22_fa19_s, lay21_fa2_c, lay21_fa1_c, lay22_fa20_s, lay22_fa20_c);
wire lay22_ha0_s, lay22_ha0_c;
half_adder lay22_ha0(lay22_fa20_s, lay21_fa0_c, lay22_ha0_s, lay22_ha0_c);
assign prod[22] = lay22_ha0_s;

wire lay23_fa0_s, lay23_fa0_c;
full_adder lay23_fa0(a23b0, a22b1, a21b2, lay23_fa0_s, lay23_fa0_c);
wire lay23_fa1_s, lay23_fa1_c;
full_adder lay23_fa1(lay23_fa0_s, a20b3, a19b4, lay23_fa1_s, lay23_fa1_c);
wire lay23_fa2_s, lay23_fa2_c;
full_adder lay23_fa2(lay23_fa1_s, a18b5, a17b6, lay23_fa2_s, lay23_fa2_c);
wire lay23_fa3_s, lay23_fa3_c;
full_adder lay23_fa3(lay23_fa2_s, a16b7, a15b8, lay23_fa3_s, lay23_fa3_c);
wire lay23_fa4_s, lay23_fa4_c;
full_adder lay23_fa4(lay23_fa3_s, a14b9, a13b10, lay23_fa4_s, lay23_fa4_c);
wire lay23_fa5_s, lay23_fa5_c;
full_adder lay23_fa5(lay23_fa4_s, a12b11, a11b12, lay23_fa5_s, lay23_fa5_c);
wire lay23_fa6_s, lay23_fa6_c;
full_adder lay23_fa6(lay23_fa5_s, a10b13, a9b14, lay23_fa6_s, lay23_fa6_c);
wire lay23_fa7_s, lay23_fa7_c;
full_adder lay23_fa7(lay23_fa6_s, a8b15, a7b16, lay23_fa7_s, lay23_fa7_c);
wire lay23_fa8_s, lay23_fa8_c;
full_adder lay23_fa8(lay23_fa7_s, a6b17, a5b18, lay23_fa8_s, lay23_fa8_c);
wire lay23_fa9_s, lay23_fa9_c;
full_adder lay23_fa9(lay23_fa8_s, a4b19, a3b20, lay23_fa9_s, lay23_fa9_c);
wire lay23_fa10_s, lay23_fa10_c;
full_adder lay23_fa10(lay23_fa9_s, a2b21, a1b22, lay23_fa10_s, lay23_fa10_c);
wire lay23_fa11_s, lay23_fa11_c;
full_adder lay23_fa11(lay23_fa10_s, a0b23, lay22_ha0_c, lay23_fa11_s, lay23_fa11_c);
wire lay23_fa12_s, lay23_fa12_c;
full_adder lay23_fa12(lay23_fa11_s, lay22_fa20_c, lay22_fa19_c, lay23_fa12_s, lay23_fa12_c);
wire lay23_fa13_s, lay23_fa13_c;
full_adder lay23_fa13(lay23_fa12_s, lay22_fa18_c, lay22_fa17_c, lay23_fa13_s, lay23_fa13_c);
wire lay23_fa14_s, lay23_fa14_c;
full_adder lay23_fa14(lay23_fa13_s, lay22_fa16_c, lay22_fa15_c, lay23_fa14_s, lay23_fa14_c);
wire lay23_fa15_s, lay23_fa15_c;
full_adder lay23_fa15(lay23_fa14_s, lay22_fa14_c, lay22_fa13_c, lay23_fa15_s, lay23_fa15_c);
wire lay23_fa16_s, lay23_fa16_c;
full_adder lay23_fa16(lay23_fa15_s, lay22_fa12_c, lay22_fa11_c, lay23_fa16_s, lay23_fa16_c);
wire lay23_fa17_s, lay23_fa17_c;
full_adder lay23_fa17(lay23_fa16_s, lay22_fa10_c, lay22_fa9_c, lay23_fa17_s, lay23_fa17_c);
wire lay23_fa18_s, lay23_fa18_c;
full_adder lay23_fa18(lay23_fa17_s, lay22_fa8_c, lay22_fa7_c, lay23_fa18_s, lay23_fa18_c);
wire lay23_fa19_s, lay23_fa19_c;
full_adder lay23_fa19(lay23_fa18_s, lay22_fa6_c, lay22_fa5_c, lay23_fa19_s, lay23_fa19_c);
wire lay23_fa20_s, lay23_fa20_c;
full_adder lay23_fa20(lay23_fa19_s, lay22_fa4_c, lay22_fa3_c, lay23_fa20_s, lay23_fa20_c);
wire lay23_fa21_s, lay23_fa21_c;
full_adder lay23_fa21(lay23_fa20_s, lay22_fa2_c, lay22_fa1_c, lay23_fa21_s, lay23_fa21_c);
wire lay23_ha0_s, lay23_ha0_c;
half_adder lay23_ha0(lay23_fa21_s, lay22_fa0_c, lay23_ha0_s, lay23_ha0_c);
assign prod[23] = lay23_ha0_s;

wire lay24_fa0_s, lay24_fa0_c;
full_adder lay24_fa0(a24b0, a23b1, a22b2, lay24_fa0_s, lay24_fa0_c);
wire lay24_fa1_s, lay24_fa1_c;
full_adder lay24_fa1(lay24_fa0_s, a21b3, a20b4, lay24_fa1_s, lay24_fa1_c);
wire lay24_fa2_s, lay24_fa2_c;
full_adder lay24_fa2(lay24_fa1_s, a19b5, a18b6, lay24_fa2_s, lay24_fa2_c);
wire lay24_fa3_s, lay24_fa3_c;
full_adder lay24_fa3(lay24_fa2_s, a17b7, a16b8, lay24_fa3_s, lay24_fa3_c);
wire lay24_fa4_s, lay24_fa4_c;
full_adder lay24_fa4(lay24_fa3_s, a15b9, a14b10, lay24_fa4_s, lay24_fa4_c);
wire lay24_fa5_s, lay24_fa5_c;
full_adder lay24_fa5(lay24_fa4_s, a13b11, a12b12, lay24_fa5_s, lay24_fa5_c);
wire lay24_fa6_s, lay24_fa6_c;
full_adder lay24_fa6(lay24_fa5_s, a11b13, a10b14, lay24_fa6_s, lay24_fa6_c);
wire lay24_fa7_s, lay24_fa7_c;
full_adder lay24_fa7(lay24_fa6_s, a9b15, a8b16, lay24_fa7_s, lay24_fa7_c);
wire lay24_fa8_s, lay24_fa8_c;
full_adder lay24_fa8(lay24_fa7_s, a7b17, a6b18, lay24_fa8_s, lay24_fa8_c);
wire lay24_fa9_s, lay24_fa9_c;
full_adder lay24_fa9(lay24_fa8_s, a5b19, a4b20, lay24_fa9_s, lay24_fa9_c);
wire lay24_fa10_s, lay24_fa10_c;
full_adder lay24_fa10(lay24_fa9_s, a3b21, a2b22, lay24_fa10_s, lay24_fa10_c);
wire lay24_fa11_s, lay24_fa11_c;
full_adder lay24_fa11(lay24_fa10_s, a1b23, a0b24, lay24_fa11_s, lay24_fa11_c);
wire lay24_fa12_s, lay24_fa12_c;
full_adder lay24_fa12(lay24_fa11_s, lay23_ha0_c, lay23_fa21_c, lay24_fa12_s, lay24_fa12_c);
wire lay24_fa13_s, lay24_fa13_c;
full_adder lay24_fa13(lay24_fa12_s, lay23_fa20_c, lay23_fa19_c, lay24_fa13_s, lay24_fa13_c);
wire lay24_fa14_s, lay24_fa14_c;
full_adder lay24_fa14(lay24_fa13_s, lay23_fa18_c, lay23_fa17_c, lay24_fa14_s, lay24_fa14_c);
wire lay24_fa15_s, lay24_fa15_c;
full_adder lay24_fa15(lay24_fa14_s, lay23_fa16_c, lay23_fa15_c, lay24_fa15_s, lay24_fa15_c);
wire lay24_fa16_s, lay24_fa16_c;
full_adder lay24_fa16(lay24_fa15_s, lay23_fa14_c, lay23_fa13_c, lay24_fa16_s, lay24_fa16_c);
wire lay24_fa17_s, lay24_fa17_c;
full_adder lay24_fa17(lay24_fa16_s, lay23_fa12_c, lay23_fa11_c, lay24_fa17_s, lay24_fa17_c);
wire lay24_fa18_s, lay24_fa18_c;
full_adder lay24_fa18(lay24_fa17_s, lay23_fa10_c, lay23_fa9_c, lay24_fa18_s, lay24_fa18_c);
wire lay24_fa19_s, lay24_fa19_c;
full_adder lay24_fa19(lay24_fa18_s, lay23_fa8_c, lay23_fa7_c, lay24_fa19_s, lay24_fa19_c);
wire lay24_fa20_s, lay24_fa20_c;
full_adder lay24_fa20(lay24_fa19_s, lay23_fa6_c, lay23_fa5_c, lay24_fa20_s, lay24_fa20_c);
wire lay24_fa21_s, lay24_fa21_c;
full_adder lay24_fa21(lay24_fa20_s, lay23_fa4_c, lay23_fa3_c, lay24_fa21_s, lay24_fa21_c);
wire lay24_fa22_s, lay24_fa22_c;
full_adder lay24_fa22(lay24_fa21_s, lay23_fa2_c, lay23_fa1_c, lay24_fa22_s, lay24_fa22_c);
wire lay24_ha0_s, lay24_ha0_c;
half_adder lay24_ha0(lay24_fa22_s, lay23_fa0_c, lay24_ha0_s, lay24_ha0_c);
assign prod[24] = lay24_ha0_s;

wire lay25_fa0_s, lay25_fa0_c;
full_adder lay25_fa0(a25b0, a24b1, a23b2, lay25_fa0_s, lay25_fa0_c);
wire lay25_fa1_s, lay25_fa1_c;
full_adder lay25_fa1(lay25_fa0_s, a22b3, a21b4, lay25_fa1_s, lay25_fa1_c);
wire lay25_fa2_s, lay25_fa2_c;
full_adder lay25_fa2(lay25_fa1_s, a20b5, a19b6, lay25_fa2_s, lay25_fa2_c);
wire lay25_fa3_s, lay25_fa3_c;
full_adder lay25_fa3(lay25_fa2_s, a18b7, a17b8, lay25_fa3_s, lay25_fa3_c);
wire lay25_fa4_s, lay25_fa4_c;
full_adder lay25_fa4(lay25_fa3_s, a16b9, a15b10, lay25_fa4_s, lay25_fa4_c);
wire lay25_fa5_s, lay25_fa5_c;
full_adder lay25_fa5(lay25_fa4_s, a14b11, a13b12, lay25_fa5_s, lay25_fa5_c);
wire lay25_fa6_s, lay25_fa6_c;
full_adder lay25_fa6(lay25_fa5_s, a12b13, a11b14, lay25_fa6_s, lay25_fa6_c);
wire lay25_fa7_s, lay25_fa7_c;
full_adder lay25_fa7(lay25_fa6_s, a10b15, a9b16, lay25_fa7_s, lay25_fa7_c);
wire lay25_fa8_s, lay25_fa8_c;
full_adder lay25_fa8(lay25_fa7_s, a8b17, a7b18, lay25_fa8_s, lay25_fa8_c);
wire lay25_fa9_s, lay25_fa9_c;
full_adder lay25_fa9(lay25_fa8_s, a6b19, a5b20, lay25_fa9_s, lay25_fa9_c);
wire lay25_fa10_s, lay25_fa10_c;
full_adder lay25_fa10(lay25_fa9_s, a4b21, a3b22, lay25_fa10_s, lay25_fa10_c);
wire lay25_fa11_s, lay25_fa11_c;
full_adder lay25_fa11(lay25_fa10_s, a2b23, a1b24, lay25_fa11_s, lay25_fa11_c);
wire lay25_fa12_s, lay25_fa12_c;
full_adder lay25_fa12(lay25_fa11_s, a0b25, lay24_ha0_c, lay25_fa12_s, lay25_fa12_c);
wire lay25_fa13_s, lay25_fa13_c;
full_adder lay25_fa13(lay25_fa12_s, lay24_fa22_c, lay24_fa21_c, lay25_fa13_s, lay25_fa13_c);
wire lay25_fa14_s, lay25_fa14_c;
full_adder lay25_fa14(lay25_fa13_s, lay24_fa20_c, lay24_fa19_c, lay25_fa14_s, lay25_fa14_c);
wire lay25_fa15_s, lay25_fa15_c;
full_adder lay25_fa15(lay25_fa14_s, lay24_fa18_c, lay24_fa17_c, lay25_fa15_s, lay25_fa15_c);
wire lay25_fa16_s, lay25_fa16_c;
full_adder lay25_fa16(lay25_fa15_s, lay24_fa16_c, lay24_fa15_c, lay25_fa16_s, lay25_fa16_c);
wire lay25_fa17_s, lay25_fa17_c;
full_adder lay25_fa17(lay25_fa16_s, lay24_fa14_c, lay24_fa13_c, lay25_fa17_s, lay25_fa17_c);
wire lay25_fa18_s, lay25_fa18_c;
full_adder lay25_fa18(lay25_fa17_s, lay24_fa12_c, lay24_fa11_c, lay25_fa18_s, lay25_fa18_c);
wire lay25_fa19_s, lay25_fa19_c;
full_adder lay25_fa19(lay25_fa18_s, lay24_fa10_c, lay24_fa9_c, lay25_fa19_s, lay25_fa19_c);
wire lay25_fa20_s, lay25_fa20_c;
full_adder lay25_fa20(lay25_fa19_s, lay24_fa8_c, lay24_fa7_c, lay25_fa20_s, lay25_fa20_c);
wire lay25_fa21_s, lay25_fa21_c;
full_adder lay25_fa21(lay25_fa20_s, lay24_fa6_c, lay24_fa5_c, lay25_fa21_s, lay25_fa21_c);
wire lay25_fa22_s, lay25_fa22_c;
full_adder lay25_fa22(lay25_fa21_s, lay24_fa4_c, lay24_fa3_c, lay25_fa22_s, lay25_fa22_c);
wire lay25_fa23_s, lay25_fa23_c;
full_adder lay25_fa23(lay25_fa22_s, lay24_fa2_c, lay24_fa1_c, lay25_fa23_s, lay25_fa23_c);
wire lay25_ha0_s, lay25_ha0_c;
half_adder lay25_ha0(lay25_fa23_s, lay24_fa0_c, lay25_ha0_s, lay25_ha0_c);
assign prod[25] = lay25_ha0_s;

wire lay26_fa0_s, lay26_fa0_c;
full_adder lay26_fa0(a26b0, a25b1, a24b2, lay26_fa0_s, lay26_fa0_c);
wire lay26_fa1_s, lay26_fa1_c;
full_adder lay26_fa1(lay26_fa0_s, a23b3, a22b4, lay26_fa1_s, lay26_fa1_c);
wire lay26_fa2_s, lay26_fa2_c;
full_adder lay26_fa2(lay26_fa1_s, a21b5, a20b6, lay26_fa2_s, lay26_fa2_c);
wire lay26_fa3_s, lay26_fa3_c;
full_adder lay26_fa3(lay26_fa2_s, a19b7, a18b8, lay26_fa3_s, lay26_fa3_c);
wire lay26_fa4_s, lay26_fa4_c;
full_adder lay26_fa4(lay26_fa3_s, a17b9, a16b10, lay26_fa4_s, lay26_fa4_c);
wire lay26_fa5_s, lay26_fa5_c;
full_adder lay26_fa5(lay26_fa4_s, a15b11, a14b12, lay26_fa5_s, lay26_fa5_c);
wire lay26_fa6_s, lay26_fa6_c;
full_adder lay26_fa6(lay26_fa5_s, a13b13, a12b14, lay26_fa6_s, lay26_fa6_c);
wire lay26_fa7_s, lay26_fa7_c;
full_adder lay26_fa7(lay26_fa6_s, a11b15, a10b16, lay26_fa7_s, lay26_fa7_c);
wire lay26_fa8_s, lay26_fa8_c;
full_adder lay26_fa8(lay26_fa7_s, a9b17, a8b18, lay26_fa8_s, lay26_fa8_c);
wire lay26_fa9_s, lay26_fa9_c;
full_adder lay26_fa9(lay26_fa8_s, a7b19, a6b20, lay26_fa9_s, lay26_fa9_c);
wire lay26_fa10_s, lay26_fa10_c;
full_adder lay26_fa10(lay26_fa9_s, a5b21, a4b22, lay26_fa10_s, lay26_fa10_c);
wire lay26_fa11_s, lay26_fa11_c;
full_adder lay26_fa11(lay26_fa10_s, a3b23, a2b24, lay26_fa11_s, lay26_fa11_c);
wire lay26_fa12_s, lay26_fa12_c;
full_adder lay26_fa12(lay26_fa11_s, a1b25, a0b26, lay26_fa12_s, lay26_fa12_c);
wire lay26_fa13_s, lay26_fa13_c;
full_adder lay26_fa13(lay26_fa12_s, lay25_ha0_c, lay25_fa23_c, lay26_fa13_s, lay26_fa13_c);
wire lay26_fa14_s, lay26_fa14_c;
full_adder lay26_fa14(lay26_fa13_s, lay25_fa22_c, lay25_fa21_c, lay26_fa14_s, lay26_fa14_c);
wire lay26_fa15_s, lay26_fa15_c;
full_adder lay26_fa15(lay26_fa14_s, lay25_fa20_c, lay25_fa19_c, lay26_fa15_s, lay26_fa15_c);
wire lay26_fa16_s, lay26_fa16_c;
full_adder lay26_fa16(lay26_fa15_s, lay25_fa18_c, lay25_fa17_c, lay26_fa16_s, lay26_fa16_c);
wire lay26_fa17_s, lay26_fa17_c;
full_adder lay26_fa17(lay26_fa16_s, lay25_fa16_c, lay25_fa15_c, lay26_fa17_s, lay26_fa17_c);
wire lay26_fa18_s, lay26_fa18_c;
full_adder lay26_fa18(lay26_fa17_s, lay25_fa14_c, lay25_fa13_c, lay26_fa18_s, lay26_fa18_c);
wire lay26_fa19_s, lay26_fa19_c;
full_adder lay26_fa19(lay26_fa18_s, lay25_fa12_c, lay25_fa11_c, lay26_fa19_s, lay26_fa19_c);
wire lay26_fa20_s, lay26_fa20_c;
full_adder lay26_fa20(lay26_fa19_s, lay25_fa10_c, lay25_fa9_c, lay26_fa20_s, lay26_fa20_c);
wire lay26_fa21_s, lay26_fa21_c;
full_adder lay26_fa21(lay26_fa20_s, lay25_fa8_c, lay25_fa7_c, lay26_fa21_s, lay26_fa21_c);
wire lay26_fa22_s, lay26_fa22_c;
full_adder lay26_fa22(lay26_fa21_s, lay25_fa6_c, lay25_fa5_c, lay26_fa22_s, lay26_fa22_c);
wire lay26_fa23_s, lay26_fa23_c;
full_adder lay26_fa23(lay26_fa22_s, lay25_fa4_c, lay25_fa3_c, lay26_fa23_s, lay26_fa23_c);
wire lay26_fa24_s, lay26_fa24_c;
full_adder lay26_fa24(lay26_fa23_s, lay25_fa2_c, lay25_fa1_c, lay26_fa24_s, lay26_fa24_c);
wire lay26_ha0_s, lay26_ha0_c;
half_adder lay26_ha0(lay26_fa24_s, lay25_fa0_c, lay26_ha0_s, lay26_ha0_c);
assign prod[26] = lay26_ha0_s;

wire lay27_fa0_s, lay27_fa0_c;
full_adder lay27_fa0(a27b0, a26b1, a25b2, lay27_fa0_s, lay27_fa0_c);
wire lay27_fa1_s, lay27_fa1_c;
full_adder lay27_fa1(lay27_fa0_s, a24b3, a23b4, lay27_fa1_s, lay27_fa1_c);
wire lay27_fa2_s, lay27_fa2_c;
full_adder lay27_fa2(lay27_fa1_s, a22b5, a21b6, lay27_fa2_s, lay27_fa2_c);
wire lay27_fa3_s, lay27_fa3_c;
full_adder lay27_fa3(lay27_fa2_s, a20b7, a19b8, lay27_fa3_s, lay27_fa3_c);
wire lay27_fa4_s, lay27_fa4_c;
full_adder lay27_fa4(lay27_fa3_s, a18b9, a17b10, lay27_fa4_s, lay27_fa4_c);
wire lay27_fa5_s, lay27_fa5_c;
full_adder lay27_fa5(lay27_fa4_s, a16b11, a15b12, lay27_fa5_s, lay27_fa5_c);
wire lay27_fa6_s, lay27_fa6_c;
full_adder lay27_fa6(lay27_fa5_s, a14b13, a13b14, lay27_fa6_s, lay27_fa6_c);
wire lay27_fa7_s, lay27_fa7_c;
full_adder lay27_fa7(lay27_fa6_s, a12b15, a11b16, lay27_fa7_s, lay27_fa7_c);
wire lay27_fa8_s, lay27_fa8_c;
full_adder lay27_fa8(lay27_fa7_s, a10b17, a9b18, lay27_fa8_s, lay27_fa8_c);
wire lay27_fa9_s, lay27_fa9_c;
full_adder lay27_fa9(lay27_fa8_s, a8b19, a7b20, lay27_fa9_s, lay27_fa9_c);
wire lay27_fa10_s, lay27_fa10_c;
full_adder lay27_fa10(lay27_fa9_s, a6b21, a5b22, lay27_fa10_s, lay27_fa10_c);
wire lay27_fa11_s, lay27_fa11_c;
full_adder lay27_fa11(lay27_fa10_s, a4b23, a3b24, lay27_fa11_s, lay27_fa11_c);
wire lay27_fa12_s, lay27_fa12_c;
full_adder lay27_fa12(lay27_fa11_s, a2b25, a1b26, lay27_fa12_s, lay27_fa12_c);
wire lay27_fa13_s, lay27_fa13_c;
full_adder lay27_fa13(lay27_fa12_s, a0b27, lay26_ha0_c, lay27_fa13_s, lay27_fa13_c);
wire lay27_fa14_s, lay27_fa14_c;
full_adder lay27_fa14(lay27_fa13_s, lay26_fa24_c, lay26_fa23_c, lay27_fa14_s, lay27_fa14_c);
wire lay27_fa15_s, lay27_fa15_c;
full_adder lay27_fa15(lay27_fa14_s, lay26_fa22_c, lay26_fa21_c, lay27_fa15_s, lay27_fa15_c);
wire lay27_fa16_s, lay27_fa16_c;
full_adder lay27_fa16(lay27_fa15_s, lay26_fa20_c, lay26_fa19_c, lay27_fa16_s, lay27_fa16_c);
wire lay27_fa17_s, lay27_fa17_c;
full_adder lay27_fa17(lay27_fa16_s, lay26_fa18_c, lay26_fa17_c, lay27_fa17_s, lay27_fa17_c);
wire lay27_fa18_s, lay27_fa18_c;
full_adder lay27_fa18(lay27_fa17_s, lay26_fa16_c, lay26_fa15_c, lay27_fa18_s, lay27_fa18_c);
wire lay27_fa19_s, lay27_fa19_c;
full_adder lay27_fa19(lay27_fa18_s, lay26_fa14_c, lay26_fa13_c, lay27_fa19_s, lay27_fa19_c);
wire lay27_fa20_s, lay27_fa20_c;
full_adder lay27_fa20(lay27_fa19_s, lay26_fa12_c, lay26_fa11_c, lay27_fa20_s, lay27_fa20_c);
wire lay27_fa21_s, lay27_fa21_c;
full_adder lay27_fa21(lay27_fa20_s, lay26_fa10_c, lay26_fa9_c, lay27_fa21_s, lay27_fa21_c);
wire lay27_fa22_s, lay27_fa22_c;
full_adder lay27_fa22(lay27_fa21_s, lay26_fa8_c, lay26_fa7_c, lay27_fa22_s, lay27_fa22_c);
wire lay27_fa23_s, lay27_fa23_c;
full_adder lay27_fa23(lay27_fa22_s, lay26_fa6_c, lay26_fa5_c, lay27_fa23_s, lay27_fa23_c);
wire lay27_fa24_s, lay27_fa24_c;
full_adder lay27_fa24(lay27_fa23_s, lay26_fa4_c, lay26_fa3_c, lay27_fa24_s, lay27_fa24_c);
wire lay27_fa25_s, lay27_fa25_c;
full_adder lay27_fa25(lay27_fa24_s, lay26_fa2_c, lay26_fa1_c, lay27_fa25_s, lay27_fa25_c);
wire lay27_ha0_s, lay27_ha0_c;
half_adder lay27_ha0(lay27_fa25_s, lay26_fa0_c, lay27_ha0_s, lay27_ha0_c);
assign prod[27] = lay27_ha0_s;

wire lay28_fa0_s, lay28_fa0_c;
full_adder lay28_fa0(a28b0, a27b1, a26b2, lay28_fa0_s, lay28_fa0_c);
wire lay28_fa1_s, lay28_fa1_c;
full_adder lay28_fa1(lay28_fa0_s, a25b3, a24b4, lay28_fa1_s, lay28_fa1_c);
wire lay28_fa2_s, lay28_fa2_c;
full_adder lay28_fa2(lay28_fa1_s, a23b5, a22b6, lay28_fa2_s, lay28_fa2_c);
wire lay28_fa3_s, lay28_fa3_c;
full_adder lay28_fa3(lay28_fa2_s, a21b7, a20b8, lay28_fa3_s, lay28_fa3_c);
wire lay28_fa4_s, lay28_fa4_c;
full_adder lay28_fa4(lay28_fa3_s, a19b9, a18b10, lay28_fa4_s, lay28_fa4_c);
wire lay28_fa5_s, lay28_fa5_c;
full_adder lay28_fa5(lay28_fa4_s, a17b11, a16b12, lay28_fa5_s, lay28_fa5_c);
wire lay28_fa6_s, lay28_fa6_c;
full_adder lay28_fa6(lay28_fa5_s, a15b13, a14b14, lay28_fa6_s, lay28_fa6_c);
wire lay28_fa7_s, lay28_fa7_c;
full_adder lay28_fa7(lay28_fa6_s, a13b15, a12b16, lay28_fa7_s, lay28_fa7_c);
wire lay28_fa8_s, lay28_fa8_c;
full_adder lay28_fa8(lay28_fa7_s, a11b17, a10b18, lay28_fa8_s, lay28_fa8_c);
wire lay28_fa9_s, lay28_fa9_c;
full_adder lay28_fa9(lay28_fa8_s, a9b19, a8b20, lay28_fa9_s, lay28_fa9_c);
wire lay28_fa10_s, lay28_fa10_c;
full_adder lay28_fa10(lay28_fa9_s, a7b21, a6b22, lay28_fa10_s, lay28_fa10_c);
wire lay28_fa11_s, lay28_fa11_c;
full_adder lay28_fa11(lay28_fa10_s, a5b23, a4b24, lay28_fa11_s, lay28_fa11_c);
wire lay28_fa12_s, lay28_fa12_c;
full_adder lay28_fa12(lay28_fa11_s, a3b25, a2b26, lay28_fa12_s, lay28_fa12_c);
wire lay28_fa13_s, lay28_fa13_c;
full_adder lay28_fa13(lay28_fa12_s, a1b27, a0b28, lay28_fa13_s, lay28_fa13_c);
wire lay28_fa14_s, lay28_fa14_c;
full_adder lay28_fa14(lay28_fa13_s, lay27_ha0_c, lay27_fa25_c, lay28_fa14_s, lay28_fa14_c);
wire lay28_fa15_s, lay28_fa15_c;
full_adder lay28_fa15(lay28_fa14_s, lay27_fa24_c, lay27_fa23_c, lay28_fa15_s, lay28_fa15_c);
wire lay28_fa16_s, lay28_fa16_c;
full_adder lay28_fa16(lay28_fa15_s, lay27_fa22_c, lay27_fa21_c, lay28_fa16_s, lay28_fa16_c);
wire lay28_fa17_s, lay28_fa17_c;
full_adder lay28_fa17(lay28_fa16_s, lay27_fa20_c, lay27_fa19_c, lay28_fa17_s, lay28_fa17_c);
wire lay28_fa18_s, lay28_fa18_c;
full_adder lay28_fa18(lay28_fa17_s, lay27_fa18_c, lay27_fa17_c, lay28_fa18_s, lay28_fa18_c);
wire lay28_fa19_s, lay28_fa19_c;
full_adder lay28_fa19(lay28_fa18_s, lay27_fa16_c, lay27_fa15_c, lay28_fa19_s, lay28_fa19_c);
wire lay28_fa20_s, lay28_fa20_c;
full_adder lay28_fa20(lay28_fa19_s, lay27_fa14_c, lay27_fa13_c, lay28_fa20_s, lay28_fa20_c);
wire lay28_fa21_s, lay28_fa21_c;
full_adder lay28_fa21(lay28_fa20_s, lay27_fa12_c, lay27_fa11_c, lay28_fa21_s, lay28_fa21_c);
wire lay28_fa22_s, lay28_fa22_c;
full_adder lay28_fa22(lay28_fa21_s, lay27_fa10_c, lay27_fa9_c, lay28_fa22_s, lay28_fa22_c);
wire lay28_fa23_s, lay28_fa23_c;
full_adder lay28_fa23(lay28_fa22_s, lay27_fa8_c, lay27_fa7_c, lay28_fa23_s, lay28_fa23_c);
wire lay28_fa24_s, lay28_fa24_c;
full_adder lay28_fa24(lay28_fa23_s, lay27_fa6_c, lay27_fa5_c, lay28_fa24_s, lay28_fa24_c);
wire lay28_fa25_s, lay28_fa25_c;
full_adder lay28_fa25(lay28_fa24_s, lay27_fa4_c, lay27_fa3_c, lay28_fa25_s, lay28_fa25_c);
wire lay28_fa26_s, lay28_fa26_c;
full_adder lay28_fa26(lay28_fa25_s, lay27_fa2_c, lay27_fa1_c, lay28_fa26_s, lay28_fa26_c);
wire lay28_ha0_s, lay28_ha0_c;
half_adder lay28_ha0(lay28_fa26_s, lay27_fa0_c, lay28_ha0_s, lay28_ha0_c);
assign prod[28] = lay28_ha0_s;

wire lay29_fa0_s, lay29_fa0_c;
full_adder lay29_fa0(a29b0, a28b1, a27b2, lay29_fa0_s, lay29_fa0_c);
wire lay29_fa1_s, lay29_fa1_c;
full_adder lay29_fa1(lay29_fa0_s, a26b3, a25b4, lay29_fa1_s, lay29_fa1_c);
wire lay29_fa2_s, lay29_fa2_c;
full_adder lay29_fa2(lay29_fa1_s, a24b5, a23b6, lay29_fa2_s, lay29_fa2_c);
wire lay29_fa3_s, lay29_fa3_c;
full_adder lay29_fa3(lay29_fa2_s, a22b7, a21b8, lay29_fa3_s, lay29_fa3_c);
wire lay29_fa4_s, lay29_fa4_c;
full_adder lay29_fa4(lay29_fa3_s, a20b9, a19b10, lay29_fa4_s, lay29_fa4_c);
wire lay29_fa5_s, lay29_fa5_c;
full_adder lay29_fa5(lay29_fa4_s, a18b11, a17b12, lay29_fa5_s, lay29_fa5_c);
wire lay29_fa6_s, lay29_fa6_c;
full_adder lay29_fa6(lay29_fa5_s, a16b13, a15b14, lay29_fa6_s, lay29_fa6_c);
wire lay29_fa7_s, lay29_fa7_c;
full_adder lay29_fa7(lay29_fa6_s, a14b15, a13b16, lay29_fa7_s, lay29_fa7_c);
wire lay29_fa8_s, lay29_fa8_c;
full_adder lay29_fa8(lay29_fa7_s, a12b17, a11b18, lay29_fa8_s, lay29_fa8_c);
wire lay29_fa9_s, lay29_fa9_c;
full_adder lay29_fa9(lay29_fa8_s, a10b19, a9b20, lay29_fa9_s, lay29_fa9_c);
wire lay29_fa10_s, lay29_fa10_c;
full_adder lay29_fa10(lay29_fa9_s, a8b21, a7b22, lay29_fa10_s, lay29_fa10_c);
wire lay29_fa11_s, lay29_fa11_c;
full_adder lay29_fa11(lay29_fa10_s, a6b23, a5b24, lay29_fa11_s, lay29_fa11_c);
wire lay29_fa12_s, lay29_fa12_c;
full_adder lay29_fa12(lay29_fa11_s, a4b25, a3b26, lay29_fa12_s, lay29_fa12_c);
wire lay29_fa13_s, lay29_fa13_c;
full_adder lay29_fa13(lay29_fa12_s, a2b27, a1b28, lay29_fa13_s, lay29_fa13_c);
wire lay29_fa14_s, lay29_fa14_c;
full_adder lay29_fa14(lay29_fa13_s, a0b29, lay28_ha0_c, lay29_fa14_s, lay29_fa14_c);
wire lay29_fa15_s, lay29_fa15_c;
full_adder lay29_fa15(lay29_fa14_s, lay28_fa26_c, lay28_fa25_c, lay29_fa15_s, lay29_fa15_c);
wire lay29_fa16_s, lay29_fa16_c;
full_adder lay29_fa16(lay29_fa15_s, lay28_fa24_c, lay28_fa23_c, lay29_fa16_s, lay29_fa16_c);
wire lay29_fa17_s, lay29_fa17_c;
full_adder lay29_fa17(lay29_fa16_s, lay28_fa22_c, lay28_fa21_c, lay29_fa17_s, lay29_fa17_c);
wire lay29_fa18_s, lay29_fa18_c;
full_adder lay29_fa18(lay29_fa17_s, lay28_fa20_c, lay28_fa19_c, lay29_fa18_s, lay29_fa18_c);
wire lay29_fa19_s, lay29_fa19_c;
full_adder lay29_fa19(lay29_fa18_s, lay28_fa18_c, lay28_fa17_c, lay29_fa19_s, lay29_fa19_c);
wire lay29_fa20_s, lay29_fa20_c;
full_adder lay29_fa20(lay29_fa19_s, lay28_fa16_c, lay28_fa15_c, lay29_fa20_s, lay29_fa20_c);
wire lay29_fa21_s, lay29_fa21_c;
full_adder lay29_fa21(lay29_fa20_s, lay28_fa14_c, lay28_fa13_c, lay29_fa21_s, lay29_fa21_c);
wire lay29_fa22_s, lay29_fa22_c;
full_adder lay29_fa22(lay29_fa21_s, lay28_fa12_c, lay28_fa11_c, lay29_fa22_s, lay29_fa22_c);
wire lay29_fa23_s, lay29_fa23_c;
full_adder lay29_fa23(lay29_fa22_s, lay28_fa10_c, lay28_fa9_c, lay29_fa23_s, lay29_fa23_c);
wire lay29_fa24_s, lay29_fa24_c;
full_adder lay29_fa24(lay29_fa23_s, lay28_fa8_c, lay28_fa7_c, lay29_fa24_s, lay29_fa24_c);
wire lay29_fa25_s, lay29_fa25_c;
full_adder lay29_fa25(lay29_fa24_s, lay28_fa6_c, lay28_fa5_c, lay29_fa25_s, lay29_fa25_c);
wire lay29_fa26_s, lay29_fa26_c;
full_adder lay29_fa26(lay29_fa25_s, lay28_fa4_c, lay28_fa3_c, lay29_fa26_s, lay29_fa26_c);
wire lay29_fa27_s, lay29_fa27_c;
full_adder lay29_fa27(lay29_fa26_s, lay28_fa2_c, lay28_fa1_c, lay29_fa27_s, lay29_fa27_c);
wire lay29_ha0_s, lay29_ha0_c;
half_adder lay29_ha0(lay29_fa27_s, lay28_fa0_c, lay29_ha0_s, lay29_ha0_c);
assign prod[29] = lay29_ha0_s;

wire lay30_fa0_s, lay30_fa0_c;
full_adder lay30_fa0(a30b0, a29b1, a28b2, lay30_fa0_s, lay30_fa0_c);
wire lay30_fa1_s, lay30_fa1_c;
full_adder lay30_fa1(lay30_fa0_s, a27b3, a26b4, lay30_fa1_s, lay30_fa1_c);
wire lay30_fa2_s, lay30_fa2_c;
full_adder lay30_fa2(lay30_fa1_s, a25b5, a24b6, lay30_fa2_s, lay30_fa2_c);
wire lay30_fa3_s, lay30_fa3_c;
full_adder lay30_fa3(lay30_fa2_s, a23b7, a22b8, lay30_fa3_s, lay30_fa3_c);
wire lay30_fa4_s, lay30_fa4_c;
full_adder lay30_fa4(lay30_fa3_s, a21b9, a20b10, lay30_fa4_s, lay30_fa4_c);
wire lay30_fa5_s, lay30_fa5_c;
full_adder lay30_fa5(lay30_fa4_s, a19b11, a18b12, lay30_fa5_s, lay30_fa5_c);
wire lay30_fa6_s, lay30_fa6_c;
full_adder lay30_fa6(lay30_fa5_s, a17b13, a16b14, lay30_fa6_s, lay30_fa6_c);
wire lay30_fa7_s, lay30_fa7_c;
full_adder lay30_fa7(lay30_fa6_s, a15b15, a14b16, lay30_fa7_s, lay30_fa7_c);
wire lay30_fa8_s, lay30_fa8_c;
full_adder lay30_fa8(lay30_fa7_s, a13b17, a12b18, lay30_fa8_s, lay30_fa8_c);
wire lay30_fa9_s, lay30_fa9_c;
full_adder lay30_fa9(lay30_fa8_s, a11b19, a10b20, lay30_fa9_s, lay30_fa9_c);
wire lay30_fa10_s, lay30_fa10_c;
full_adder lay30_fa10(lay30_fa9_s, a9b21, a8b22, lay30_fa10_s, lay30_fa10_c);
wire lay30_fa11_s, lay30_fa11_c;
full_adder lay30_fa11(lay30_fa10_s, a7b23, a6b24, lay30_fa11_s, lay30_fa11_c);
wire lay30_fa12_s, lay30_fa12_c;
full_adder lay30_fa12(lay30_fa11_s, a5b25, a4b26, lay30_fa12_s, lay30_fa12_c);
wire lay30_fa13_s, lay30_fa13_c;
full_adder lay30_fa13(lay30_fa12_s, a3b27, a2b28, lay30_fa13_s, lay30_fa13_c);
wire lay30_fa14_s, lay30_fa14_c;
full_adder lay30_fa14(lay30_fa13_s, a1b29, a0b30, lay30_fa14_s, lay30_fa14_c);
wire lay30_fa15_s, lay30_fa15_c;
full_adder lay30_fa15(lay30_fa14_s, lay29_ha0_c, lay29_fa27_c, lay30_fa15_s, lay30_fa15_c);
wire lay30_fa16_s, lay30_fa16_c;
full_adder lay30_fa16(lay30_fa15_s, lay29_fa26_c, lay29_fa25_c, lay30_fa16_s, lay30_fa16_c);
wire lay30_fa17_s, lay30_fa17_c;
full_adder lay30_fa17(lay30_fa16_s, lay29_fa24_c, lay29_fa23_c, lay30_fa17_s, lay30_fa17_c);
wire lay30_fa18_s, lay30_fa18_c;
full_adder lay30_fa18(lay30_fa17_s, lay29_fa22_c, lay29_fa21_c, lay30_fa18_s, lay30_fa18_c);
wire lay30_fa19_s, lay30_fa19_c;
full_adder lay30_fa19(lay30_fa18_s, lay29_fa20_c, lay29_fa19_c, lay30_fa19_s, lay30_fa19_c);
wire lay30_fa20_s, lay30_fa20_c;
full_adder lay30_fa20(lay30_fa19_s, lay29_fa18_c, lay29_fa17_c, lay30_fa20_s, lay30_fa20_c);
wire lay30_fa21_s, lay30_fa21_c;
full_adder lay30_fa21(lay30_fa20_s, lay29_fa16_c, lay29_fa15_c, lay30_fa21_s, lay30_fa21_c);
wire lay30_fa22_s, lay30_fa22_c;
full_adder lay30_fa22(lay30_fa21_s, lay29_fa14_c, lay29_fa13_c, lay30_fa22_s, lay30_fa22_c);
wire lay30_fa23_s, lay30_fa23_c;
full_adder lay30_fa23(lay30_fa22_s, lay29_fa12_c, lay29_fa11_c, lay30_fa23_s, lay30_fa23_c);
wire lay30_fa24_s, lay30_fa24_c;
full_adder lay30_fa24(lay30_fa23_s, lay29_fa10_c, lay29_fa9_c, lay30_fa24_s, lay30_fa24_c);
wire lay30_fa25_s, lay30_fa25_c;
full_adder lay30_fa25(lay30_fa24_s, lay29_fa8_c, lay29_fa7_c, lay30_fa25_s, lay30_fa25_c);
wire lay30_fa26_s, lay30_fa26_c;
full_adder lay30_fa26(lay30_fa25_s, lay29_fa6_c, lay29_fa5_c, lay30_fa26_s, lay30_fa26_c);
wire lay30_fa27_s, lay30_fa27_c;
full_adder lay30_fa27(lay30_fa26_s, lay29_fa4_c, lay29_fa3_c, lay30_fa27_s, lay30_fa27_c);
wire lay30_fa28_s, lay30_fa28_c;
full_adder lay30_fa28(lay30_fa27_s, lay29_fa2_c, lay29_fa1_c, lay30_fa28_s, lay30_fa28_c);
wire lay30_ha0_s, lay30_ha0_c;
half_adder lay30_ha0(lay30_fa28_s, lay29_fa0_c, lay30_ha0_s, lay30_ha0_c);
assign prod[30] = lay30_ha0_s;

wire lay31_fa0_s, lay31_fa0_c;
full_adder lay31_fa0(a31b0, a30b1, a29b2, lay31_fa0_s, lay31_fa0_c);
wire lay31_fa1_s, lay31_fa1_c;
full_adder lay31_fa1(lay31_fa0_s, a28b3, a27b4, lay31_fa1_s, lay31_fa1_c);
wire lay31_fa2_s, lay31_fa2_c;
full_adder lay31_fa2(lay31_fa1_s, a26b5, a25b6, lay31_fa2_s, lay31_fa2_c);
wire lay31_fa3_s, lay31_fa3_c;
full_adder lay31_fa3(lay31_fa2_s, a24b7, a23b8, lay31_fa3_s, lay31_fa3_c);
wire lay31_fa4_s, lay31_fa4_c;
full_adder lay31_fa4(lay31_fa3_s, a22b9, a21b10, lay31_fa4_s, lay31_fa4_c);
wire lay31_fa5_s, lay31_fa5_c;
full_adder lay31_fa5(lay31_fa4_s, a20b11, a19b12, lay31_fa5_s, lay31_fa5_c);
wire lay31_fa6_s, lay31_fa6_c;
full_adder lay31_fa6(lay31_fa5_s, a18b13, a17b14, lay31_fa6_s, lay31_fa6_c);
wire lay31_fa7_s, lay31_fa7_c;
full_adder lay31_fa7(lay31_fa6_s, a16b15, a15b16, lay31_fa7_s, lay31_fa7_c);
wire lay31_fa8_s, lay31_fa8_c;
full_adder lay31_fa8(lay31_fa7_s, a14b17, a13b18, lay31_fa8_s, lay31_fa8_c);
wire lay31_fa9_s, lay31_fa9_c;
full_adder lay31_fa9(lay31_fa8_s, a12b19, a11b20, lay31_fa9_s, lay31_fa9_c);
wire lay31_fa10_s, lay31_fa10_c;
full_adder lay31_fa10(lay31_fa9_s, a10b21, a9b22, lay31_fa10_s, lay31_fa10_c);
wire lay31_fa11_s, lay31_fa11_c;
full_adder lay31_fa11(lay31_fa10_s, a8b23, a7b24, lay31_fa11_s, lay31_fa11_c);
wire lay31_fa12_s, lay31_fa12_c;
full_adder lay31_fa12(lay31_fa11_s, a6b25, a5b26, lay31_fa12_s, lay31_fa12_c);
wire lay31_fa13_s, lay31_fa13_c;
full_adder lay31_fa13(lay31_fa12_s, a4b27, a3b28, lay31_fa13_s, lay31_fa13_c);
wire lay31_fa14_s, lay31_fa14_c;
full_adder lay31_fa14(lay31_fa13_s, a2b29, a1b30, lay31_fa14_s, lay31_fa14_c);
wire lay31_fa15_s, lay31_fa15_c;
full_adder lay31_fa15(lay31_fa14_s, a0b31, lay30_ha0_c, lay31_fa15_s, lay31_fa15_c);
wire lay31_fa16_s, lay31_fa16_c;
full_adder lay31_fa16(lay31_fa15_s, lay30_fa28_c, lay30_fa27_c, lay31_fa16_s, lay31_fa16_c);
wire lay31_fa17_s, lay31_fa17_c;
full_adder lay31_fa17(lay31_fa16_s, lay30_fa26_c, lay30_fa25_c, lay31_fa17_s, lay31_fa17_c);
wire lay31_fa18_s, lay31_fa18_c;
full_adder lay31_fa18(lay31_fa17_s, lay30_fa24_c, lay30_fa23_c, lay31_fa18_s, lay31_fa18_c);
wire lay31_fa19_s, lay31_fa19_c;
full_adder lay31_fa19(lay31_fa18_s, lay30_fa22_c, lay30_fa21_c, lay31_fa19_s, lay31_fa19_c);
wire lay31_fa20_s, lay31_fa20_c;
full_adder lay31_fa20(lay31_fa19_s, lay30_fa20_c, lay30_fa19_c, lay31_fa20_s, lay31_fa20_c);
wire lay31_fa21_s, lay31_fa21_c;
full_adder lay31_fa21(lay31_fa20_s, lay30_fa18_c, lay30_fa17_c, lay31_fa21_s, lay31_fa21_c);
wire lay31_fa22_s, lay31_fa22_c;
full_adder lay31_fa22(lay31_fa21_s, lay30_fa16_c, lay30_fa15_c, lay31_fa22_s, lay31_fa22_c);
wire lay31_fa23_s, lay31_fa23_c;
full_adder lay31_fa23(lay31_fa22_s, lay30_fa14_c, lay30_fa13_c, lay31_fa23_s, lay31_fa23_c);
wire lay31_fa24_s, lay31_fa24_c;
full_adder lay31_fa24(lay31_fa23_s, lay30_fa12_c, lay30_fa11_c, lay31_fa24_s, lay31_fa24_c);
wire lay31_fa25_s, lay31_fa25_c;
full_adder lay31_fa25(lay31_fa24_s, lay30_fa10_c, lay30_fa9_c, lay31_fa25_s, lay31_fa25_c);
wire lay31_fa26_s, lay31_fa26_c;
full_adder lay31_fa26(lay31_fa25_s, lay30_fa8_c, lay30_fa7_c, lay31_fa26_s, lay31_fa26_c);
wire lay31_fa27_s, lay31_fa27_c;
full_adder lay31_fa27(lay31_fa26_s, lay30_fa6_c, lay30_fa5_c, lay31_fa27_s, lay31_fa27_c);
wire lay31_fa28_s, lay31_fa28_c;
full_adder lay31_fa28(lay31_fa27_s, lay30_fa4_c, lay30_fa3_c, lay31_fa28_s, lay31_fa28_c);
wire lay31_fa29_s, lay31_fa29_c;
full_adder lay31_fa29(lay31_fa28_s, lay30_fa2_c, lay30_fa1_c, lay31_fa29_s, lay31_fa29_c);
wire lay31_ha0_s, lay31_ha0_c;
half_adder lay31_ha0(lay31_fa29_s, lay30_fa0_c, lay31_ha0_s, lay31_ha0_c);
assign prod[31] = lay31_ha0_s;

wire lay32_fa0_s, lay32_fa0_c;
full_adder lay32_fa0(1'b1, a31b1, a30b2, lay32_fa0_s, lay32_fa0_c);
wire lay32_fa1_s, lay32_fa1_c;
full_adder lay32_fa1(lay32_fa0_s, a29b3, a28b4, lay32_fa1_s, lay32_fa1_c);
wire lay32_fa2_s, lay32_fa2_c;
full_adder lay32_fa2(lay32_fa1_s, a27b5, a26b6, lay32_fa2_s, lay32_fa2_c);
wire lay32_fa3_s, lay32_fa3_c;
full_adder lay32_fa3(lay32_fa2_s, a25b7, a24b8, lay32_fa3_s, lay32_fa3_c);
wire lay32_fa4_s, lay32_fa4_c;
full_adder lay32_fa4(lay32_fa3_s, a23b9, a22b10, lay32_fa4_s, lay32_fa4_c);
wire lay32_fa5_s, lay32_fa5_c;
full_adder lay32_fa5(lay32_fa4_s, a21b11, a20b12, lay32_fa5_s, lay32_fa5_c);
wire lay32_fa6_s, lay32_fa6_c;
full_adder lay32_fa6(lay32_fa5_s, a19b13, a18b14, lay32_fa6_s, lay32_fa6_c);
wire lay32_fa7_s, lay32_fa7_c;
full_adder lay32_fa7(lay32_fa6_s, a17b15, a16b16, lay32_fa7_s, lay32_fa7_c);
wire lay32_fa8_s, lay32_fa8_c;
full_adder lay32_fa8(lay32_fa7_s, a15b17, a14b18, lay32_fa8_s, lay32_fa8_c);
wire lay32_fa9_s, lay32_fa9_c;
full_adder lay32_fa9(lay32_fa8_s, a13b19, a12b20, lay32_fa9_s, lay32_fa9_c);
wire lay32_fa10_s, lay32_fa10_c;
full_adder lay32_fa10(lay32_fa9_s, a11b21, a10b22, lay32_fa10_s, lay32_fa10_c);
wire lay32_fa11_s, lay32_fa11_c;
full_adder lay32_fa11(lay32_fa10_s, a9b23, a8b24, lay32_fa11_s, lay32_fa11_c);
wire lay32_fa12_s, lay32_fa12_c;
full_adder lay32_fa12(lay32_fa11_s, a7b25, a6b26, lay32_fa12_s, lay32_fa12_c);
wire lay32_fa13_s, lay32_fa13_c;
full_adder lay32_fa13(lay32_fa12_s, a5b27, a4b28, lay32_fa13_s, lay32_fa13_c);
wire lay32_fa14_s, lay32_fa14_c;
full_adder lay32_fa14(lay32_fa13_s, a3b29, a2b30, lay32_fa14_s, lay32_fa14_c);
wire lay32_fa15_s, lay32_fa15_c;
full_adder lay32_fa15(lay32_fa14_s, a1b31, lay31_ha0_c, lay32_fa15_s, lay32_fa15_c);
wire lay32_fa16_s, lay32_fa16_c;
full_adder lay32_fa16(lay32_fa15_s, lay31_fa29_c, lay31_fa28_c, lay32_fa16_s, lay32_fa16_c);
wire lay32_fa17_s, lay32_fa17_c;
full_adder lay32_fa17(lay32_fa16_s, lay31_fa27_c, lay31_fa26_c, lay32_fa17_s, lay32_fa17_c);
wire lay32_fa18_s, lay32_fa18_c;
full_adder lay32_fa18(lay32_fa17_s, lay31_fa25_c, lay31_fa24_c, lay32_fa18_s, lay32_fa18_c);
wire lay32_fa19_s, lay32_fa19_c;
full_adder lay32_fa19(lay32_fa18_s, lay31_fa23_c, lay31_fa22_c, lay32_fa19_s, lay32_fa19_c);
wire lay32_fa20_s, lay32_fa20_c;
full_adder lay32_fa20(lay32_fa19_s, lay31_fa21_c, lay31_fa20_c, lay32_fa20_s, lay32_fa20_c);
wire lay32_fa21_s, lay32_fa21_c;
full_adder lay32_fa21(lay32_fa20_s, lay31_fa19_c, lay31_fa18_c, lay32_fa21_s, lay32_fa21_c);
wire lay32_fa22_s, lay32_fa22_c;
full_adder lay32_fa22(lay32_fa21_s, lay31_fa17_c, lay31_fa16_c, lay32_fa22_s, lay32_fa22_c);
wire lay32_fa23_s, lay32_fa23_c;
full_adder lay32_fa23(lay32_fa22_s, lay31_fa15_c, lay31_fa14_c, lay32_fa23_s, lay32_fa23_c);
wire lay32_fa24_s, lay32_fa24_c;
full_adder lay32_fa24(lay32_fa23_s, lay31_fa13_c, lay31_fa12_c, lay32_fa24_s, lay32_fa24_c);
wire lay32_fa25_s, lay32_fa25_c;
full_adder lay32_fa25(lay32_fa24_s, lay31_fa11_c, lay31_fa10_c, lay32_fa25_s, lay32_fa25_c);
wire lay32_fa26_s, lay32_fa26_c;
full_adder lay32_fa26(lay32_fa25_s, lay31_fa9_c, lay31_fa8_c, lay32_fa26_s, lay32_fa26_c);
wire lay32_fa27_s, lay32_fa27_c;
full_adder lay32_fa27(lay32_fa26_s, lay31_fa7_c, lay31_fa6_c, lay32_fa27_s, lay32_fa27_c);
wire lay32_fa28_s, lay32_fa28_c;
full_adder lay32_fa28(lay32_fa27_s, lay31_fa5_c, lay31_fa4_c, lay32_fa28_s, lay32_fa28_c);
wire lay32_fa29_s, lay32_fa29_c;
full_adder lay32_fa29(lay32_fa28_s, lay31_fa3_c, lay31_fa2_c, lay32_fa29_s, lay32_fa29_c);
wire lay32_fa30_s, lay32_fa30_c;
full_adder lay32_fa30(lay32_fa29_s, lay31_fa1_c, lay31_fa0_c, lay32_fa30_s, lay32_fa30_c);
assign prod[32] = lay32_fa30_s;

wire lay33_fa0_s, lay33_fa0_c;
full_adder lay33_fa0(a31b2, a30b3, a29b4, lay33_fa0_s, lay33_fa0_c);
wire lay33_fa1_s, lay33_fa1_c;
full_adder lay33_fa1(lay33_fa0_s, a28b5, a27b6, lay33_fa1_s, lay33_fa1_c);
wire lay33_fa2_s, lay33_fa2_c;
full_adder lay33_fa2(lay33_fa1_s, a26b7, a25b8, lay33_fa2_s, lay33_fa2_c);
wire lay33_fa3_s, lay33_fa3_c;
full_adder lay33_fa3(lay33_fa2_s, a24b9, a23b10, lay33_fa3_s, lay33_fa3_c);
wire lay33_fa4_s, lay33_fa4_c;
full_adder lay33_fa4(lay33_fa3_s, a22b11, a21b12, lay33_fa4_s, lay33_fa4_c);
wire lay33_fa5_s, lay33_fa5_c;
full_adder lay33_fa5(lay33_fa4_s, a20b13, a19b14, lay33_fa5_s, lay33_fa5_c);
wire lay33_fa6_s, lay33_fa6_c;
full_adder lay33_fa6(lay33_fa5_s, a18b15, a17b16, lay33_fa6_s, lay33_fa6_c);
wire lay33_fa7_s, lay33_fa7_c;
full_adder lay33_fa7(lay33_fa6_s, a16b17, a15b18, lay33_fa7_s, lay33_fa7_c);
wire lay33_fa8_s, lay33_fa8_c;
full_adder lay33_fa8(lay33_fa7_s, a14b19, a13b20, lay33_fa8_s, lay33_fa8_c);
wire lay33_fa9_s, lay33_fa9_c;
full_adder lay33_fa9(lay33_fa8_s, a12b21, a11b22, lay33_fa9_s, lay33_fa9_c);
wire lay33_fa10_s, lay33_fa10_c;
full_adder lay33_fa10(lay33_fa9_s, a10b23, a9b24, lay33_fa10_s, lay33_fa10_c);
wire lay33_fa11_s, lay33_fa11_c;
full_adder lay33_fa11(lay33_fa10_s, a8b25, a7b26, lay33_fa11_s, lay33_fa11_c);
wire lay33_fa12_s, lay33_fa12_c;
full_adder lay33_fa12(lay33_fa11_s, a6b27, a5b28, lay33_fa12_s, lay33_fa12_c);
wire lay33_fa13_s, lay33_fa13_c;
full_adder lay33_fa13(lay33_fa12_s, a4b29, a3b30, lay33_fa13_s, lay33_fa13_c);
wire lay33_fa14_s, lay33_fa14_c;
full_adder lay33_fa14(lay33_fa13_s, a2b31, lay32_fa30_c, lay33_fa14_s, lay33_fa14_c);
wire lay33_fa15_s, lay33_fa15_c;
full_adder lay33_fa15(lay33_fa14_s, lay32_fa29_c, lay32_fa28_c, lay33_fa15_s, lay33_fa15_c);
wire lay33_fa16_s, lay33_fa16_c;
full_adder lay33_fa16(lay33_fa15_s, lay32_fa27_c, lay32_fa26_c, lay33_fa16_s, lay33_fa16_c);
wire lay33_fa17_s, lay33_fa17_c;
full_adder lay33_fa17(lay33_fa16_s, lay32_fa25_c, lay32_fa24_c, lay33_fa17_s, lay33_fa17_c);
wire lay33_fa18_s, lay33_fa18_c;
full_adder lay33_fa18(lay33_fa17_s, lay32_fa23_c, lay32_fa22_c, lay33_fa18_s, lay33_fa18_c);
wire lay33_fa19_s, lay33_fa19_c;
full_adder lay33_fa19(lay33_fa18_s, lay32_fa21_c, lay32_fa20_c, lay33_fa19_s, lay33_fa19_c);
wire lay33_fa20_s, lay33_fa20_c;
full_adder lay33_fa20(lay33_fa19_s, lay32_fa19_c, lay32_fa18_c, lay33_fa20_s, lay33_fa20_c);
wire lay33_fa21_s, lay33_fa21_c;
full_adder lay33_fa21(lay33_fa20_s, lay32_fa17_c, lay32_fa16_c, lay33_fa21_s, lay33_fa21_c);
wire lay33_fa22_s, lay33_fa22_c;
full_adder lay33_fa22(lay33_fa21_s, lay32_fa15_c, lay32_fa14_c, lay33_fa22_s, lay33_fa22_c);
wire lay33_fa23_s, lay33_fa23_c;
full_adder lay33_fa23(lay33_fa22_s, lay32_fa13_c, lay32_fa12_c, lay33_fa23_s, lay33_fa23_c);
wire lay33_fa24_s, lay33_fa24_c;
full_adder lay33_fa24(lay33_fa23_s, lay32_fa11_c, lay32_fa10_c, lay33_fa24_s, lay33_fa24_c);
wire lay33_fa25_s, lay33_fa25_c;
full_adder lay33_fa25(lay33_fa24_s, lay32_fa9_c, lay32_fa8_c, lay33_fa25_s, lay33_fa25_c);
wire lay33_fa26_s, lay33_fa26_c;
full_adder lay33_fa26(lay33_fa25_s, lay32_fa7_c, lay32_fa6_c, lay33_fa26_s, lay33_fa26_c);
wire lay33_fa27_s, lay33_fa27_c;
full_adder lay33_fa27(lay33_fa26_s, lay32_fa5_c, lay32_fa4_c, lay33_fa27_s, lay33_fa27_c);
wire lay33_fa28_s, lay33_fa28_c;
full_adder lay33_fa28(lay33_fa27_s, lay32_fa3_c, lay32_fa2_c, lay33_fa28_s, lay33_fa28_c);
wire lay33_fa29_s, lay33_fa29_c;
full_adder lay33_fa29(lay33_fa28_s, lay32_fa1_c, lay32_fa0_c, lay33_fa29_s, lay33_fa29_c);
assign prod[33] = lay33_fa29_s;

wire lay34_fa0_s, lay34_fa0_c;
full_adder lay34_fa0(a31b3, a30b4, a29b5, lay34_fa0_s, lay34_fa0_c);
wire lay34_fa1_s, lay34_fa1_c;
full_adder lay34_fa1(lay34_fa0_s, a28b6, a27b7, lay34_fa1_s, lay34_fa1_c);
wire lay34_fa2_s, lay34_fa2_c;
full_adder lay34_fa2(lay34_fa1_s, a26b8, a25b9, lay34_fa2_s, lay34_fa2_c);
wire lay34_fa3_s, lay34_fa3_c;
full_adder lay34_fa3(lay34_fa2_s, a24b10, a23b11, lay34_fa3_s, lay34_fa3_c);
wire lay34_fa4_s, lay34_fa4_c;
full_adder lay34_fa4(lay34_fa3_s, a22b12, a21b13, lay34_fa4_s, lay34_fa4_c);
wire lay34_fa5_s, lay34_fa5_c;
full_adder lay34_fa5(lay34_fa4_s, a20b14, a19b15, lay34_fa5_s, lay34_fa5_c);
wire lay34_fa6_s, lay34_fa6_c;
full_adder lay34_fa6(lay34_fa5_s, a18b16, a17b17, lay34_fa6_s, lay34_fa6_c);
wire lay34_fa7_s, lay34_fa7_c;
full_adder lay34_fa7(lay34_fa6_s, a16b18, a15b19, lay34_fa7_s, lay34_fa7_c);
wire lay34_fa8_s, lay34_fa8_c;
full_adder lay34_fa8(lay34_fa7_s, a14b20, a13b21, lay34_fa8_s, lay34_fa8_c);
wire lay34_fa9_s, lay34_fa9_c;
full_adder lay34_fa9(lay34_fa8_s, a12b22, a11b23, lay34_fa9_s, lay34_fa9_c);
wire lay34_fa10_s, lay34_fa10_c;
full_adder lay34_fa10(lay34_fa9_s, a10b24, a9b25, lay34_fa10_s, lay34_fa10_c);
wire lay34_fa11_s, lay34_fa11_c;
full_adder lay34_fa11(lay34_fa10_s, a8b26, a7b27, lay34_fa11_s, lay34_fa11_c);
wire lay34_fa12_s, lay34_fa12_c;
full_adder lay34_fa12(lay34_fa11_s, a6b28, a5b29, lay34_fa12_s, lay34_fa12_c);
wire lay34_fa13_s, lay34_fa13_c;
full_adder lay34_fa13(lay34_fa12_s, a4b30, a3b31, lay34_fa13_s, lay34_fa13_c);
wire lay34_fa14_s, lay34_fa14_c;
full_adder lay34_fa14(lay34_fa13_s, lay33_fa29_c, lay33_fa28_c, lay34_fa14_s, lay34_fa14_c);
wire lay34_fa15_s, lay34_fa15_c;
full_adder lay34_fa15(lay34_fa14_s, lay33_fa27_c, lay33_fa26_c, lay34_fa15_s, lay34_fa15_c);
wire lay34_fa16_s, lay34_fa16_c;
full_adder lay34_fa16(lay34_fa15_s, lay33_fa25_c, lay33_fa24_c, lay34_fa16_s, lay34_fa16_c);
wire lay34_fa17_s, lay34_fa17_c;
full_adder lay34_fa17(lay34_fa16_s, lay33_fa23_c, lay33_fa22_c, lay34_fa17_s, lay34_fa17_c);
wire lay34_fa18_s, lay34_fa18_c;
full_adder lay34_fa18(lay34_fa17_s, lay33_fa21_c, lay33_fa20_c, lay34_fa18_s, lay34_fa18_c);
wire lay34_fa19_s, lay34_fa19_c;
full_adder lay34_fa19(lay34_fa18_s, lay33_fa19_c, lay33_fa18_c, lay34_fa19_s, lay34_fa19_c);
wire lay34_fa20_s, lay34_fa20_c;
full_adder lay34_fa20(lay34_fa19_s, lay33_fa17_c, lay33_fa16_c, lay34_fa20_s, lay34_fa20_c);
wire lay34_fa21_s, lay34_fa21_c;
full_adder lay34_fa21(lay34_fa20_s, lay33_fa15_c, lay33_fa14_c, lay34_fa21_s, lay34_fa21_c);
wire lay34_fa22_s, lay34_fa22_c;
full_adder lay34_fa22(lay34_fa21_s, lay33_fa13_c, lay33_fa12_c, lay34_fa22_s, lay34_fa22_c);
wire lay34_fa23_s, lay34_fa23_c;
full_adder lay34_fa23(lay34_fa22_s, lay33_fa11_c, lay33_fa10_c, lay34_fa23_s, lay34_fa23_c);
wire lay34_fa24_s, lay34_fa24_c;
full_adder lay34_fa24(lay34_fa23_s, lay33_fa9_c, lay33_fa8_c, lay34_fa24_s, lay34_fa24_c);
wire lay34_fa25_s, lay34_fa25_c;
full_adder lay34_fa25(lay34_fa24_s, lay33_fa7_c, lay33_fa6_c, lay34_fa25_s, lay34_fa25_c);
wire lay34_fa26_s, lay34_fa26_c;
full_adder lay34_fa26(lay34_fa25_s, lay33_fa5_c, lay33_fa4_c, lay34_fa26_s, lay34_fa26_c);
wire lay34_fa27_s, lay34_fa27_c;
full_adder lay34_fa27(lay34_fa26_s, lay33_fa3_c, lay33_fa2_c, lay34_fa27_s, lay34_fa27_c);
wire lay34_fa28_s, lay34_fa28_c;
full_adder lay34_fa28(lay34_fa27_s, lay33_fa1_c, lay33_fa0_c, lay34_fa28_s, lay34_fa28_c);
assign prod[34] = lay34_fa28_s;

wire lay35_fa0_s, lay35_fa0_c;
full_adder lay35_fa0(a31b4, a30b5, a29b6, lay35_fa0_s, lay35_fa0_c);
wire lay35_fa1_s, lay35_fa1_c;
full_adder lay35_fa1(lay35_fa0_s, a28b7, a27b8, lay35_fa1_s, lay35_fa1_c);
wire lay35_fa2_s, lay35_fa2_c;
full_adder lay35_fa2(lay35_fa1_s, a26b9, a25b10, lay35_fa2_s, lay35_fa2_c);
wire lay35_fa3_s, lay35_fa3_c;
full_adder lay35_fa3(lay35_fa2_s, a24b11, a23b12, lay35_fa3_s, lay35_fa3_c);
wire lay35_fa4_s, lay35_fa4_c;
full_adder lay35_fa4(lay35_fa3_s, a22b13, a21b14, lay35_fa4_s, lay35_fa4_c);
wire lay35_fa5_s, lay35_fa5_c;
full_adder lay35_fa5(lay35_fa4_s, a20b15, a19b16, lay35_fa5_s, lay35_fa5_c);
wire lay35_fa6_s, lay35_fa6_c;
full_adder lay35_fa6(lay35_fa5_s, a18b17, a17b18, lay35_fa6_s, lay35_fa6_c);
wire lay35_fa7_s, lay35_fa7_c;
full_adder lay35_fa7(lay35_fa6_s, a16b19, a15b20, lay35_fa7_s, lay35_fa7_c);
wire lay35_fa8_s, lay35_fa8_c;
full_adder lay35_fa8(lay35_fa7_s, a14b21, a13b22, lay35_fa8_s, lay35_fa8_c);
wire lay35_fa9_s, lay35_fa9_c;
full_adder lay35_fa9(lay35_fa8_s, a12b23, a11b24, lay35_fa9_s, lay35_fa9_c);
wire lay35_fa10_s, lay35_fa10_c;
full_adder lay35_fa10(lay35_fa9_s, a10b25, a9b26, lay35_fa10_s, lay35_fa10_c);
wire lay35_fa11_s, lay35_fa11_c;
full_adder lay35_fa11(lay35_fa10_s, a8b27, a7b28, lay35_fa11_s, lay35_fa11_c);
wire lay35_fa12_s, lay35_fa12_c;
full_adder lay35_fa12(lay35_fa11_s, a6b29, a5b30, lay35_fa12_s, lay35_fa12_c);
wire lay35_fa13_s, lay35_fa13_c;
full_adder lay35_fa13(lay35_fa12_s, a4b31, lay34_fa28_c, lay35_fa13_s, lay35_fa13_c);
wire lay35_fa14_s, lay35_fa14_c;
full_adder lay35_fa14(lay35_fa13_s, lay34_fa27_c, lay34_fa26_c, lay35_fa14_s, lay35_fa14_c);
wire lay35_fa15_s, lay35_fa15_c;
full_adder lay35_fa15(lay35_fa14_s, lay34_fa25_c, lay34_fa24_c, lay35_fa15_s, lay35_fa15_c);
wire lay35_fa16_s, lay35_fa16_c;
full_adder lay35_fa16(lay35_fa15_s, lay34_fa23_c, lay34_fa22_c, lay35_fa16_s, lay35_fa16_c);
wire lay35_fa17_s, lay35_fa17_c;
full_adder lay35_fa17(lay35_fa16_s, lay34_fa21_c, lay34_fa20_c, lay35_fa17_s, lay35_fa17_c);
wire lay35_fa18_s, lay35_fa18_c;
full_adder lay35_fa18(lay35_fa17_s, lay34_fa19_c, lay34_fa18_c, lay35_fa18_s, lay35_fa18_c);
wire lay35_fa19_s, lay35_fa19_c;
full_adder lay35_fa19(lay35_fa18_s, lay34_fa17_c, lay34_fa16_c, lay35_fa19_s, lay35_fa19_c);
wire lay35_fa20_s, lay35_fa20_c;
full_adder lay35_fa20(lay35_fa19_s, lay34_fa15_c, lay34_fa14_c, lay35_fa20_s, lay35_fa20_c);
wire lay35_fa21_s, lay35_fa21_c;
full_adder lay35_fa21(lay35_fa20_s, lay34_fa13_c, lay34_fa12_c, lay35_fa21_s, lay35_fa21_c);
wire lay35_fa22_s, lay35_fa22_c;
full_adder lay35_fa22(lay35_fa21_s, lay34_fa11_c, lay34_fa10_c, lay35_fa22_s, lay35_fa22_c);
wire lay35_fa23_s, lay35_fa23_c;
full_adder lay35_fa23(lay35_fa22_s, lay34_fa9_c, lay34_fa8_c, lay35_fa23_s, lay35_fa23_c);
wire lay35_fa24_s, lay35_fa24_c;
full_adder lay35_fa24(lay35_fa23_s, lay34_fa7_c, lay34_fa6_c, lay35_fa24_s, lay35_fa24_c);
wire lay35_fa25_s, lay35_fa25_c;
full_adder lay35_fa25(lay35_fa24_s, lay34_fa5_c, lay34_fa4_c, lay35_fa25_s, lay35_fa25_c);
wire lay35_fa26_s, lay35_fa26_c;
full_adder lay35_fa26(lay35_fa25_s, lay34_fa3_c, lay34_fa2_c, lay35_fa26_s, lay35_fa26_c);
wire lay35_fa27_s, lay35_fa27_c;
full_adder lay35_fa27(lay35_fa26_s, lay34_fa1_c, lay34_fa0_c, lay35_fa27_s, lay35_fa27_c);
assign prod[35] = lay35_fa27_s;

wire lay36_fa0_s, lay36_fa0_c;
full_adder lay36_fa0(a31b5, a30b6, a29b7, lay36_fa0_s, lay36_fa0_c);
wire lay36_fa1_s, lay36_fa1_c;
full_adder lay36_fa1(lay36_fa0_s, a28b8, a27b9, lay36_fa1_s, lay36_fa1_c);
wire lay36_fa2_s, lay36_fa2_c;
full_adder lay36_fa2(lay36_fa1_s, a26b10, a25b11, lay36_fa2_s, lay36_fa2_c);
wire lay36_fa3_s, lay36_fa3_c;
full_adder lay36_fa3(lay36_fa2_s, a24b12, a23b13, lay36_fa3_s, lay36_fa3_c);
wire lay36_fa4_s, lay36_fa4_c;
full_adder lay36_fa4(lay36_fa3_s, a22b14, a21b15, lay36_fa4_s, lay36_fa4_c);
wire lay36_fa5_s, lay36_fa5_c;
full_adder lay36_fa5(lay36_fa4_s, a20b16, a19b17, lay36_fa5_s, lay36_fa5_c);
wire lay36_fa6_s, lay36_fa6_c;
full_adder lay36_fa6(lay36_fa5_s, a18b18, a17b19, lay36_fa6_s, lay36_fa6_c);
wire lay36_fa7_s, lay36_fa7_c;
full_adder lay36_fa7(lay36_fa6_s, a16b20, a15b21, lay36_fa7_s, lay36_fa7_c);
wire lay36_fa8_s, lay36_fa8_c;
full_adder lay36_fa8(lay36_fa7_s, a14b22, a13b23, lay36_fa8_s, lay36_fa8_c);
wire lay36_fa9_s, lay36_fa9_c;
full_adder lay36_fa9(lay36_fa8_s, a12b24, a11b25, lay36_fa9_s, lay36_fa9_c);
wire lay36_fa10_s, lay36_fa10_c;
full_adder lay36_fa10(lay36_fa9_s, a10b26, a9b27, lay36_fa10_s, lay36_fa10_c);
wire lay36_fa11_s, lay36_fa11_c;
full_adder lay36_fa11(lay36_fa10_s, a8b28, a7b29, lay36_fa11_s, lay36_fa11_c);
wire lay36_fa12_s, lay36_fa12_c;
full_adder lay36_fa12(lay36_fa11_s, a6b30, a5b31, lay36_fa12_s, lay36_fa12_c);
wire lay36_fa13_s, lay36_fa13_c;
full_adder lay36_fa13(lay36_fa12_s, lay35_fa27_c, lay35_fa26_c, lay36_fa13_s, lay36_fa13_c);
wire lay36_fa14_s, lay36_fa14_c;
full_adder lay36_fa14(lay36_fa13_s, lay35_fa25_c, lay35_fa24_c, lay36_fa14_s, lay36_fa14_c);
wire lay36_fa15_s, lay36_fa15_c;
full_adder lay36_fa15(lay36_fa14_s, lay35_fa23_c, lay35_fa22_c, lay36_fa15_s, lay36_fa15_c);
wire lay36_fa16_s, lay36_fa16_c;
full_adder lay36_fa16(lay36_fa15_s, lay35_fa21_c, lay35_fa20_c, lay36_fa16_s, lay36_fa16_c);
wire lay36_fa17_s, lay36_fa17_c;
full_adder lay36_fa17(lay36_fa16_s, lay35_fa19_c, lay35_fa18_c, lay36_fa17_s, lay36_fa17_c);
wire lay36_fa18_s, lay36_fa18_c;
full_adder lay36_fa18(lay36_fa17_s, lay35_fa17_c, lay35_fa16_c, lay36_fa18_s, lay36_fa18_c);
wire lay36_fa19_s, lay36_fa19_c;
full_adder lay36_fa19(lay36_fa18_s, lay35_fa15_c, lay35_fa14_c, lay36_fa19_s, lay36_fa19_c);
wire lay36_fa20_s, lay36_fa20_c;
full_adder lay36_fa20(lay36_fa19_s, lay35_fa13_c, lay35_fa12_c, lay36_fa20_s, lay36_fa20_c);
wire lay36_fa21_s, lay36_fa21_c;
full_adder lay36_fa21(lay36_fa20_s, lay35_fa11_c, lay35_fa10_c, lay36_fa21_s, lay36_fa21_c);
wire lay36_fa22_s, lay36_fa22_c;
full_adder lay36_fa22(lay36_fa21_s, lay35_fa9_c, lay35_fa8_c, lay36_fa22_s, lay36_fa22_c);
wire lay36_fa23_s, lay36_fa23_c;
full_adder lay36_fa23(lay36_fa22_s, lay35_fa7_c, lay35_fa6_c, lay36_fa23_s, lay36_fa23_c);
wire lay36_fa24_s, lay36_fa24_c;
full_adder lay36_fa24(lay36_fa23_s, lay35_fa5_c, lay35_fa4_c, lay36_fa24_s, lay36_fa24_c);
wire lay36_fa25_s, lay36_fa25_c;
full_adder lay36_fa25(lay36_fa24_s, lay35_fa3_c, lay35_fa2_c, lay36_fa25_s, lay36_fa25_c);
wire lay36_fa26_s, lay36_fa26_c;
full_adder lay36_fa26(lay36_fa25_s, lay35_fa1_c, lay35_fa0_c, lay36_fa26_s, lay36_fa26_c);
assign prod[36] = lay36_fa26_s;

wire lay37_fa0_s, lay37_fa0_c;
full_adder lay37_fa0(a31b6, a30b7, a29b8, lay37_fa0_s, lay37_fa0_c);
wire lay37_fa1_s, lay37_fa1_c;
full_adder lay37_fa1(lay37_fa0_s, a28b9, a27b10, lay37_fa1_s, lay37_fa1_c);
wire lay37_fa2_s, lay37_fa2_c;
full_adder lay37_fa2(lay37_fa1_s, a26b11, a25b12, lay37_fa2_s, lay37_fa2_c);
wire lay37_fa3_s, lay37_fa3_c;
full_adder lay37_fa3(lay37_fa2_s, a24b13, a23b14, lay37_fa3_s, lay37_fa3_c);
wire lay37_fa4_s, lay37_fa4_c;
full_adder lay37_fa4(lay37_fa3_s, a22b15, a21b16, lay37_fa4_s, lay37_fa4_c);
wire lay37_fa5_s, lay37_fa5_c;
full_adder lay37_fa5(lay37_fa4_s, a20b17, a19b18, lay37_fa5_s, lay37_fa5_c);
wire lay37_fa6_s, lay37_fa6_c;
full_adder lay37_fa6(lay37_fa5_s, a18b19, a17b20, lay37_fa6_s, lay37_fa6_c);
wire lay37_fa7_s, lay37_fa7_c;
full_adder lay37_fa7(lay37_fa6_s, a16b21, a15b22, lay37_fa7_s, lay37_fa7_c);
wire lay37_fa8_s, lay37_fa8_c;
full_adder lay37_fa8(lay37_fa7_s, a14b23, a13b24, lay37_fa8_s, lay37_fa8_c);
wire lay37_fa9_s, lay37_fa9_c;
full_adder lay37_fa9(lay37_fa8_s, a12b25, a11b26, lay37_fa9_s, lay37_fa9_c);
wire lay37_fa10_s, lay37_fa10_c;
full_adder lay37_fa10(lay37_fa9_s, a10b27, a9b28, lay37_fa10_s, lay37_fa10_c);
wire lay37_fa11_s, lay37_fa11_c;
full_adder lay37_fa11(lay37_fa10_s, a8b29, a7b30, lay37_fa11_s, lay37_fa11_c);
wire lay37_fa12_s, lay37_fa12_c;
full_adder lay37_fa12(lay37_fa11_s, a6b31, lay36_fa26_c, lay37_fa12_s, lay37_fa12_c);
wire lay37_fa13_s, lay37_fa13_c;
full_adder lay37_fa13(lay37_fa12_s, lay36_fa25_c, lay36_fa24_c, lay37_fa13_s, lay37_fa13_c);
wire lay37_fa14_s, lay37_fa14_c;
full_adder lay37_fa14(lay37_fa13_s, lay36_fa23_c, lay36_fa22_c, lay37_fa14_s, lay37_fa14_c);
wire lay37_fa15_s, lay37_fa15_c;
full_adder lay37_fa15(lay37_fa14_s, lay36_fa21_c, lay36_fa20_c, lay37_fa15_s, lay37_fa15_c);
wire lay37_fa16_s, lay37_fa16_c;
full_adder lay37_fa16(lay37_fa15_s, lay36_fa19_c, lay36_fa18_c, lay37_fa16_s, lay37_fa16_c);
wire lay37_fa17_s, lay37_fa17_c;
full_adder lay37_fa17(lay37_fa16_s, lay36_fa17_c, lay36_fa16_c, lay37_fa17_s, lay37_fa17_c);
wire lay37_fa18_s, lay37_fa18_c;
full_adder lay37_fa18(lay37_fa17_s, lay36_fa15_c, lay36_fa14_c, lay37_fa18_s, lay37_fa18_c);
wire lay37_fa19_s, lay37_fa19_c;
full_adder lay37_fa19(lay37_fa18_s, lay36_fa13_c, lay36_fa12_c, lay37_fa19_s, lay37_fa19_c);
wire lay37_fa20_s, lay37_fa20_c;
full_adder lay37_fa20(lay37_fa19_s, lay36_fa11_c, lay36_fa10_c, lay37_fa20_s, lay37_fa20_c);
wire lay37_fa21_s, lay37_fa21_c;
full_adder lay37_fa21(lay37_fa20_s, lay36_fa9_c, lay36_fa8_c, lay37_fa21_s, lay37_fa21_c);
wire lay37_fa22_s, lay37_fa22_c;
full_adder lay37_fa22(lay37_fa21_s, lay36_fa7_c, lay36_fa6_c, lay37_fa22_s, lay37_fa22_c);
wire lay37_fa23_s, lay37_fa23_c;
full_adder lay37_fa23(lay37_fa22_s, lay36_fa5_c, lay36_fa4_c, lay37_fa23_s, lay37_fa23_c);
wire lay37_fa24_s, lay37_fa24_c;
full_adder lay37_fa24(lay37_fa23_s, lay36_fa3_c, lay36_fa2_c, lay37_fa24_s, lay37_fa24_c);
wire lay37_fa25_s, lay37_fa25_c;
full_adder lay37_fa25(lay37_fa24_s, lay36_fa1_c, lay36_fa0_c, lay37_fa25_s, lay37_fa25_c);
assign prod[37] = lay37_fa25_s;

wire lay38_fa0_s, lay38_fa0_c;
full_adder lay38_fa0(a31b7, a30b8, a29b9, lay38_fa0_s, lay38_fa0_c);
wire lay38_fa1_s, lay38_fa1_c;
full_adder lay38_fa1(lay38_fa0_s, a28b10, a27b11, lay38_fa1_s, lay38_fa1_c);
wire lay38_fa2_s, lay38_fa2_c;
full_adder lay38_fa2(lay38_fa1_s, a26b12, a25b13, lay38_fa2_s, lay38_fa2_c);
wire lay38_fa3_s, lay38_fa3_c;
full_adder lay38_fa3(lay38_fa2_s, a24b14, a23b15, lay38_fa3_s, lay38_fa3_c);
wire lay38_fa4_s, lay38_fa4_c;
full_adder lay38_fa4(lay38_fa3_s, a22b16, a21b17, lay38_fa4_s, lay38_fa4_c);
wire lay38_fa5_s, lay38_fa5_c;
full_adder lay38_fa5(lay38_fa4_s, a20b18, a19b19, lay38_fa5_s, lay38_fa5_c);
wire lay38_fa6_s, lay38_fa6_c;
full_adder lay38_fa6(lay38_fa5_s, a18b20, a17b21, lay38_fa6_s, lay38_fa6_c);
wire lay38_fa7_s, lay38_fa7_c;
full_adder lay38_fa7(lay38_fa6_s, a16b22, a15b23, lay38_fa7_s, lay38_fa7_c);
wire lay38_fa8_s, lay38_fa8_c;
full_adder lay38_fa8(lay38_fa7_s, a14b24, a13b25, lay38_fa8_s, lay38_fa8_c);
wire lay38_fa9_s, lay38_fa9_c;
full_adder lay38_fa9(lay38_fa8_s, a12b26, a11b27, lay38_fa9_s, lay38_fa9_c);
wire lay38_fa10_s, lay38_fa10_c;
full_adder lay38_fa10(lay38_fa9_s, a10b28, a9b29, lay38_fa10_s, lay38_fa10_c);
wire lay38_fa11_s, lay38_fa11_c;
full_adder lay38_fa11(lay38_fa10_s, a8b30, a7b31, lay38_fa11_s, lay38_fa11_c);
wire lay38_fa12_s, lay38_fa12_c;
full_adder lay38_fa12(lay38_fa11_s, lay37_fa25_c, lay37_fa24_c, lay38_fa12_s, lay38_fa12_c);
wire lay38_fa13_s, lay38_fa13_c;
full_adder lay38_fa13(lay38_fa12_s, lay37_fa23_c, lay37_fa22_c, lay38_fa13_s, lay38_fa13_c);
wire lay38_fa14_s, lay38_fa14_c;
full_adder lay38_fa14(lay38_fa13_s, lay37_fa21_c, lay37_fa20_c, lay38_fa14_s, lay38_fa14_c);
wire lay38_fa15_s, lay38_fa15_c;
full_adder lay38_fa15(lay38_fa14_s, lay37_fa19_c, lay37_fa18_c, lay38_fa15_s, lay38_fa15_c);
wire lay38_fa16_s, lay38_fa16_c;
full_adder lay38_fa16(lay38_fa15_s, lay37_fa17_c, lay37_fa16_c, lay38_fa16_s, lay38_fa16_c);
wire lay38_fa17_s, lay38_fa17_c;
full_adder lay38_fa17(lay38_fa16_s, lay37_fa15_c, lay37_fa14_c, lay38_fa17_s, lay38_fa17_c);
wire lay38_fa18_s, lay38_fa18_c;
full_adder lay38_fa18(lay38_fa17_s, lay37_fa13_c, lay37_fa12_c, lay38_fa18_s, lay38_fa18_c);
wire lay38_fa19_s, lay38_fa19_c;
full_adder lay38_fa19(lay38_fa18_s, lay37_fa11_c, lay37_fa10_c, lay38_fa19_s, lay38_fa19_c);
wire lay38_fa20_s, lay38_fa20_c;
full_adder lay38_fa20(lay38_fa19_s, lay37_fa9_c, lay37_fa8_c, lay38_fa20_s, lay38_fa20_c);
wire lay38_fa21_s, lay38_fa21_c;
full_adder lay38_fa21(lay38_fa20_s, lay37_fa7_c, lay37_fa6_c, lay38_fa21_s, lay38_fa21_c);
wire lay38_fa22_s, lay38_fa22_c;
full_adder lay38_fa22(lay38_fa21_s, lay37_fa5_c, lay37_fa4_c, lay38_fa22_s, lay38_fa22_c);
wire lay38_fa23_s, lay38_fa23_c;
full_adder lay38_fa23(lay38_fa22_s, lay37_fa3_c, lay37_fa2_c, lay38_fa23_s, lay38_fa23_c);
wire lay38_fa24_s, lay38_fa24_c;
full_adder lay38_fa24(lay38_fa23_s, lay37_fa1_c, lay37_fa0_c, lay38_fa24_s, lay38_fa24_c);
assign prod[38] = lay38_fa24_s;

wire lay39_fa0_s, lay39_fa0_c;
full_adder lay39_fa0(a31b8, a30b9, a29b10, lay39_fa0_s, lay39_fa0_c);
wire lay39_fa1_s, lay39_fa1_c;
full_adder lay39_fa1(lay39_fa0_s, a28b11, a27b12, lay39_fa1_s, lay39_fa1_c);
wire lay39_fa2_s, lay39_fa2_c;
full_adder lay39_fa2(lay39_fa1_s, a26b13, a25b14, lay39_fa2_s, lay39_fa2_c);
wire lay39_fa3_s, lay39_fa3_c;
full_adder lay39_fa3(lay39_fa2_s, a24b15, a23b16, lay39_fa3_s, lay39_fa3_c);
wire lay39_fa4_s, lay39_fa4_c;
full_adder lay39_fa4(lay39_fa3_s, a22b17, a21b18, lay39_fa4_s, lay39_fa4_c);
wire lay39_fa5_s, lay39_fa5_c;
full_adder lay39_fa5(lay39_fa4_s, a20b19, a19b20, lay39_fa5_s, lay39_fa5_c);
wire lay39_fa6_s, lay39_fa6_c;
full_adder lay39_fa6(lay39_fa5_s, a18b21, a17b22, lay39_fa6_s, lay39_fa6_c);
wire lay39_fa7_s, lay39_fa7_c;
full_adder lay39_fa7(lay39_fa6_s, a16b23, a15b24, lay39_fa7_s, lay39_fa7_c);
wire lay39_fa8_s, lay39_fa8_c;
full_adder lay39_fa8(lay39_fa7_s, a14b25, a13b26, lay39_fa8_s, lay39_fa8_c);
wire lay39_fa9_s, lay39_fa9_c;
full_adder lay39_fa9(lay39_fa8_s, a12b27, a11b28, lay39_fa9_s, lay39_fa9_c);
wire lay39_fa10_s, lay39_fa10_c;
full_adder lay39_fa10(lay39_fa9_s, a10b29, a9b30, lay39_fa10_s, lay39_fa10_c);
wire lay39_fa11_s, lay39_fa11_c;
full_adder lay39_fa11(lay39_fa10_s, a8b31, lay38_fa24_c, lay39_fa11_s, lay39_fa11_c);
wire lay39_fa12_s, lay39_fa12_c;
full_adder lay39_fa12(lay39_fa11_s, lay38_fa23_c, lay38_fa22_c, lay39_fa12_s, lay39_fa12_c);
wire lay39_fa13_s, lay39_fa13_c;
full_adder lay39_fa13(lay39_fa12_s, lay38_fa21_c, lay38_fa20_c, lay39_fa13_s, lay39_fa13_c);
wire lay39_fa14_s, lay39_fa14_c;
full_adder lay39_fa14(lay39_fa13_s, lay38_fa19_c, lay38_fa18_c, lay39_fa14_s, lay39_fa14_c);
wire lay39_fa15_s, lay39_fa15_c;
full_adder lay39_fa15(lay39_fa14_s, lay38_fa17_c, lay38_fa16_c, lay39_fa15_s, lay39_fa15_c);
wire lay39_fa16_s, lay39_fa16_c;
full_adder lay39_fa16(lay39_fa15_s, lay38_fa15_c, lay38_fa14_c, lay39_fa16_s, lay39_fa16_c);
wire lay39_fa17_s, lay39_fa17_c;
full_adder lay39_fa17(lay39_fa16_s, lay38_fa13_c, lay38_fa12_c, lay39_fa17_s, lay39_fa17_c);
wire lay39_fa18_s, lay39_fa18_c;
full_adder lay39_fa18(lay39_fa17_s, lay38_fa11_c, lay38_fa10_c, lay39_fa18_s, lay39_fa18_c);
wire lay39_fa19_s, lay39_fa19_c;
full_adder lay39_fa19(lay39_fa18_s, lay38_fa9_c, lay38_fa8_c, lay39_fa19_s, lay39_fa19_c);
wire lay39_fa20_s, lay39_fa20_c;
full_adder lay39_fa20(lay39_fa19_s, lay38_fa7_c, lay38_fa6_c, lay39_fa20_s, lay39_fa20_c);
wire lay39_fa21_s, lay39_fa21_c;
full_adder lay39_fa21(lay39_fa20_s, lay38_fa5_c, lay38_fa4_c, lay39_fa21_s, lay39_fa21_c);
wire lay39_fa22_s, lay39_fa22_c;
full_adder lay39_fa22(lay39_fa21_s, lay38_fa3_c, lay38_fa2_c, lay39_fa22_s, lay39_fa22_c);
wire lay39_fa23_s, lay39_fa23_c;
full_adder lay39_fa23(lay39_fa22_s, lay38_fa1_c, lay38_fa0_c, lay39_fa23_s, lay39_fa23_c);
assign prod[39] = lay39_fa23_s;

wire lay40_fa0_s, lay40_fa0_c;
full_adder lay40_fa0(a31b9, a30b10, a29b11, lay40_fa0_s, lay40_fa0_c);
wire lay40_fa1_s, lay40_fa1_c;
full_adder lay40_fa1(lay40_fa0_s, a28b12, a27b13, lay40_fa1_s, lay40_fa1_c);
wire lay40_fa2_s, lay40_fa2_c;
full_adder lay40_fa2(lay40_fa1_s, a26b14, a25b15, lay40_fa2_s, lay40_fa2_c);
wire lay40_fa3_s, lay40_fa3_c;
full_adder lay40_fa3(lay40_fa2_s, a24b16, a23b17, lay40_fa3_s, lay40_fa3_c);
wire lay40_fa4_s, lay40_fa4_c;
full_adder lay40_fa4(lay40_fa3_s, a22b18, a21b19, lay40_fa4_s, lay40_fa4_c);
wire lay40_fa5_s, lay40_fa5_c;
full_adder lay40_fa5(lay40_fa4_s, a20b20, a19b21, lay40_fa5_s, lay40_fa5_c);
wire lay40_fa6_s, lay40_fa6_c;
full_adder lay40_fa6(lay40_fa5_s, a18b22, a17b23, lay40_fa6_s, lay40_fa6_c);
wire lay40_fa7_s, lay40_fa7_c;
full_adder lay40_fa7(lay40_fa6_s, a16b24, a15b25, lay40_fa7_s, lay40_fa7_c);
wire lay40_fa8_s, lay40_fa8_c;
full_adder lay40_fa8(lay40_fa7_s, a14b26, a13b27, lay40_fa8_s, lay40_fa8_c);
wire lay40_fa9_s, lay40_fa9_c;
full_adder lay40_fa9(lay40_fa8_s, a12b28, a11b29, lay40_fa9_s, lay40_fa9_c);
wire lay40_fa10_s, lay40_fa10_c;
full_adder lay40_fa10(lay40_fa9_s, a10b30, a9b31, lay40_fa10_s, lay40_fa10_c);
wire lay40_fa11_s, lay40_fa11_c;
full_adder lay40_fa11(lay40_fa10_s, lay39_fa23_c, lay39_fa22_c, lay40_fa11_s, lay40_fa11_c);
wire lay40_fa12_s, lay40_fa12_c;
full_adder lay40_fa12(lay40_fa11_s, lay39_fa21_c, lay39_fa20_c, lay40_fa12_s, lay40_fa12_c);
wire lay40_fa13_s, lay40_fa13_c;
full_adder lay40_fa13(lay40_fa12_s, lay39_fa19_c, lay39_fa18_c, lay40_fa13_s, lay40_fa13_c);
wire lay40_fa14_s, lay40_fa14_c;
full_adder lay40_fa14(lay40_fa13_s, lay39_fa17_c, lay39_fa16_c, lay40_fa14_s, lay40_fa14_c);
wire lay40_fa15_s, lay40_fa15_c;
full_adder lay40_fa15(lay40_fa14_s, lay39_fa15_c, lay39_fa14_c, lay40_fa15_s, lay40_fa15_c);
wire lay40_fa16_s, lay40_fa16_c;
full_adder lay40_fa16(lay40_fa15_s, lay39_fa13_c, lay39_fa12_c, lay40_fa16_s, lay40_fa16_c);
wire lay40_fa17_s, lay40_fa17_c;
full_adder lay40_fa17(lay40_fa16_s, lay39_fa11_c, lay39_fa10_c, lay40_fa17_s, lay40_fa17_c);
wire lay40_fa18_s, lay40_fa18_c;
full_adder lay40_fa18(lay40_fa17_s, lay39_fa9_c, lay39_fa8_c, lay40_fa18_s, lay40_fa18_c);
wire lay40_fa19_s, lay40_fa19_c;
full_adder lay40_fa19(lay40_fa18_s, lay39_fa7_c, lay39_fa6_c, lay40_fa19_s, lay40_fa19_c);
wire lay40_fa20_s, lay40_fa20_c;
full_adder lay40_fa20(lay40_fa19_s, lay39_fa5_c, lay39_fa4_c, lay40_fa20_s, lay40_fa20_c);
wire lay40_fa21_s, lay40_fa21_c;
full_adder lay40_fa21(lay40_fa20_s, lay39_fa3_c, lay39_fa2_c, lay40_fa21_s, lay40_fa21_c);
wire lay40_fa22_s, lay40_fa22_c;
full_adder lay40_fa22(lay40_fa21_s, lay39_fa1_c, lay39_fa0_c, lay40_fa22_s, lay40_fa22_c);
assign prod[40] = lay40_fa22_s;

wire lay41_fa0_s, lay41_fa0_c;
full_adder lay41_fa0(a31b10, a30b11, a29b12, lay41_fa0_s, lay41_fa0_c);
wire lay41_fa1_s, lay41_fa1_c;
full_adder lay41_fa1(lay41_fa0_s, a28b13, a27b14, lay41_fa1_s, lay41_fa1_c);
wire lay41_fa2_s, lay41_fa2_c;
full_adder lay41_fa2(lay41_fa1_s, a26b15, a25b16, lay41_fa2_s, lay41_fa2_c);
wire lay41_fa3_s, lay41_fa3_c;
full_adder lay41_fa3(lay41_fa2_s, a24b17, a23b18, lay41_fa3_s, lay41_fa3_c);
wire lay41_fa4_s, lay41_fa4_c;
full_adder lay41_fa4(lay41_fa3_s, a22b19, a21b20, lay41_fa4_s, lay41_fa4_c);
wire lay41_fa5_s, lay41_fa5_c;
full_adder lay41_fa5(lay41_fa4_s, a20b21, a19b22, lay41_fa5_s, lay41_fa5_c);
wire lay41_fa6_s, lay41_fa6_c;
full_adder lay41_fa6(lay41_fa5_s, a18b23, a17b24, lay41_fa6_s, lay41_fa6_c);
wire lay41_fa7_s, lay41_fa7_c;
full_adder lay41_fa7(lay41_fa6_s, a16b25, a15b26, lay41_fa7_s, lay41_fa7_c);
wire lay41_fa8_s, lay41_fa8_c;
full_adder lay41_fa8(lay41_fa7_s, a14b27, a13b28, lay41_fa8_s, lay41_fa8_c);
wire lay41_fa9_s, lay41_fa9_c;
full_adder lay41_fa9(lay41_fa8_s, a12b29, a11b30, lay41_fa9_s, lay41_fa9_c);
wire lay41_fa10_s, lay41_fa10_c;
full_adder lay41_fa10(lay41_fa9_s, a10b31, lay40_fa22_c, lay41_fa10_s, lay41_fa10_c);
wire lay41_fa11_s, lay41_fa11_c;
full_adder lay41_fa11(lay41_fa10_s, lay40_fa21_c, lay40_fa20_c, lay41_fa11_s, lay41_fa11_c);
wire lay41_fa12_s, lay41_fa12_c;
full_adder lay41_fa12(lay41_fa11_s, lay40_fa19_c, lay40_fa18_c, lay41_fa12_s, lay41_fa12_c);
wire lay41_fa13_s, lay41_fa13_c;
full_adder lay41_fa13(lay41_fa12_s, lay40_fa17_c, lay40_fa16_c, lay41_fa13_s, lay41_fa13_c);
wire lay41_fa14_s, lay41_fa14_c;
full_adder lay41_fa14(lay41_fa13_s, lay40_fa15_c, lay40_fa14_c, lay41_fa14_s, lay41_fa14_c);
wire lay41_fa15_s, lay41_fa15_c;
full_adder lay41_fa15(lay41_fa14_s, lay40_fa13_c, lay40_fa12_c, lay41_fa15_s, lay41_fa15_c);
wire lay41_fa16_s, lay41_fa16_c;
full_adder lay41_fa16(lay41_fa15_s, lay40_fa11_c, lay40_fa10_c, lay41_fa16_s, lay41_fa16_c);
wire lay41_fa17_s, lay41_fa17_c;
full_adder lay41_fa17(lay41_fa16_s, lay40_fa9_c, lay40_fa8_c, lay41_fa17_s, lay41_fa17_c);
wire lay41_fa18_s, lay41_fa18_c;
full_adder lay41_fa18(lay41_fa17_s, lay40_fa7_c, lay40_fa6_c, lay41_fa18_s, lay41_fa18_c);
wire lay41_fa19_s, lay41_fa19_c;
full_adder lay41_fa19(lay41_fa18_s, lay40_fa5_c, lay40_fa4_c, lay41_fa19_s, lay41_fa19_c);
wire lay41_fa20_s, lay41_fa20_c;
full_adder lay41_fa20(lay41_fa19_s, lay40_fa3_c, lay40_fa2_c, lay41_fa20_s, lay41_fa20_c);
wire lay41_fa21_s, lay41_fa21_c;
full_adder lay41_fa21(lay41_fa20_s, lay40_fa1_c, lay40_fa0_c, lay41_fa21_s, lay41_fa21_c);
assign prod[41] = lay41_fa21_s;

wire lay42_fa0_s, lay42_fa0_c;
full_adder lay42_fa0(a31b11, a30b12, a29b13, lay42_fa0_s, lay42_fa0_c);
wire lay42_fa1_s, lay42_fa1_c;
full_adder lay42_fa1(lay42_fa0_s, a28b14, a27b15, lay42_fa1_s, lay42_fa1_c);
wire lay42_fa2_s, lay42_fa2_c;
full_adder lay42_fa2(lay42_fa1_s, a26b16, a25b17, lay42_fa2_s, lay42_fa2_c);
wire lay42_fa3_s, lay42_fa3_c;
full_adder lay42_fa3(lay42_fa2_s, a24b18, a23b19, lay42_fa3_s, lay42_fa3_c);
wire lay42_fa4_s, lay42_fa4_c;
full_adder lay42_fa4(lay42_fa3_s, a22b20, a21b21, lay42_fa4_s, lay42_fa4_c);
wire lay42_fa5_s, lay42_fa5_c;
full_adder lay42_fa5(lay42_fa4_s, a20b22, a19b23, lay42_fa5_s, lay42_fa5_c);
wire lay42_fa6_s, lay42_fa6_c;
full_adder lay42_fa6(lay42_fa5_s, a18b24, a17b25, lay42_fa6_s, lay42_fa6_c);
wire lay42_fa7_s, lay42_fa7_c;
full_adder lay42_fa7(lay42_fa6_s, a16b26, a15b27, lay42_fa7_s, lay42_fa7_c);
wire lay42_fa8_s, lay42_fa8_c;
full_adder lay42_fa8(lay42_fa7_s, a14b28, a13b29, lay42_fa8_s, lay42_fa8_c);
wire lay42_fa9_s, lay42_fa9_c;
full_adder lay42_fa9(lay42_fa8_s, a12b30, a11b31, lay42_fa9_s, lay42_fa9_c);
wire lay42_fa10_s, lay42_fa10_c;
full_adder lay42_fa10(lay42_fa9_s, lay41_fa21_c, lay41_fa20_c, lay42_fa10_s, lay42_fa10_c);
wire lay42_fa11_s, lay42_fa11_c;
full_adder lay42_fa11(lay42_fa10_s, lay41_fa19_c, lay41_fa18_c, lay42_fa11_s, lay42_fa11_c);
wire lay42_fa12_s, lay42_fa12_c;
full_adder lay42_fa12(lay42_fa11_s, lay41_fa17_c, lay41_fa16_c, lay42_fa12_s, lay42_fa12_c);
wire lay42_fa13_s, lay42_fa13_c;
full_adder lay42_fa13(lay42_fa12_s, lay41_fa15_c, lay41_fa14_c, lay42_fa13_s, lay42_fa13_c);
wire lay42_fa14_s, lay42_fa14_c;
full_adder lay42_fa14(lay42_fa13_s, lay41_fa13_c, lay41_fa12_c, lay42_fa14_s, lay42_fa14_c);
wire lay42_fa15_s, lay42_fa15_c;
full_adder lay42_fa15(lay42_fa14_s, lay41_fa11_c, lay41_fa10_c, lay42_fa15_s, lay42_fa15_c);
wire lay42_fa16_s, lay42_fa16_c;
full_adder lay42_fa16(lay42_fa15_s, lay41_fa9_c, lay41_fa8_c, lay42_fa16_s, lay42_fa16_c);
wire lay42_fa17_s, lay42_fa17_c;
full_adder lay42_fa17(lay42_fa16_s, lay41_fa7_c, lay41_fa6_c, lay42_fa17_s, lay42_fa17_c);
wire lay42_fa18_s, lay42_fa18_c;
full_adder lay42_fa18(lay42_fa17_s, lay41_fa5_c, lay41_fa4_c, lay42_fa18_s, lay42_fa18_c);
wire lay42_fa19_s, lay42_fa19_c;
full_adder lay42_fa19(lay42_fa18_s, lay41_fa3_c, lay41_fa2_c, lay42_fa19_s, lay42_fa19_c);
wire lay42_fa20_s, lay42_fa20_c;
full_adder lay42_fa20(lay42_fa19_s, lay41_fa1_c, lay41_fa0_c, lay42_fa20_s, lay42_fa20_c);
assign prod[42] = lay42_fa20_s;

wire lay43_fa0_s, lay43_fa0_c;
full_adder lay43_fa0(a31b12, a30b13, a29b14, lay43_fa0_s, lay43_fa0_c);
wire lay43_fa1_s, lay43_fa1_c;
full_adder lay43_fa1(lay43_fa0_s, a28b15, a27b16, lay43_fa1_s, lay43_fa1_c);
wire lay43_fa2_s, lay43_fa2_c;
full_adder lay43_fa2(lay43_fa1_s, a26b17, a25b18, lay43_fa2_s, lay43_fa2_c);
wire lay43_fa3_s, lay43_fa3_c;
full_adder lay43_fa3(lay43_fa2_s, a24b19, a23b20, lay43_fa3_s, lay43_fa3_c);
wire lay43_fa4_s, lay43_fa4_c;
full_adder lay43_fa4(lay43_fa3_s, a22b21, a21b22, lay43_fa4_s, lay43_fa4_c);
wire lay43_fa5_s, lay43_fa5_c;
full_adder lay43_fa5(lay43_fa4_s, a20b23, a19b24, lay43_fa5_s, lay43_fa5_c);
wire lay43_fa6_s, lay43_fa6_c;
full_adder lay43_fa6(lay43_fa5_s, a18b25, a17b26, lay43_fa6_s, lay43_fa6_c);
wire lay43_fa7_s, lay43_fa7_c;
full_adder lay43_fa7(lay43_fa6_s, a16b27, a15b28, lay43_fa7_s, lay43_fa7_c);
wire lay43_fa8_s, lay43_fa8_c;
full_adder lay43_fa8(lay43_fa7_s, a14b29, a13b30, lay43_fa8_s, lay43_fa8_c);
wire lay43_fa9_s, lay43_fa9_c;
full_adder lay43_fa9(lay43_fa8_s, a12b31, lay42_fa20_c, lay43_fa9_s, lay43_fa9_c);
wire lay43_fa10_s, lay43_fa10_c;
full_adder lay43_fa10(lay43_fa9_s, lay42_fa19_c, lay42_fa18_c, lay43_fa10_s, lay43_fa10_c);
wire lay43_fa11_s, lay43_fa11_c;
full_adder lay43_fa11(lay43_fa10_s, lay42_fa17_c, lay42_fa16_c, lay43_fa11_s, lay43_fa11_c);
wire lay43_fa12_s, lay43_fa12_c;
full_adder lay43_fa12(lay43_fa11_s, lay42_fa15_c, lay42_fa14_c, lay43_fa12_s, lay43_fa12_c);
wire lay43_fa13_s, lay43_fa13_c;
full_adder lay43_fa13(lay43_fa12_s, lay42_fa13_c, lay42_fa12_c, lay43_fa13_s, lay43_fa13_c);
wire lay43_fa14_s, lay43_fa14_c;
full_adder lay43_fa14(lay43_fa13_s, lay42_fa11_c, lay42_fa10_c, lay43_fa14_s, lay43_fa14_c);
wire lay43_fa15_s, lay43_fa15_c;
full_adder lay43_fa15(lay43_fa14_s, lay42_fa9_c, lay42_fa8_c, lay43_fa15_s, lay43_fa15_c);
wire lay43_fa16_s, lay43_fa16_c;
full_adder lay43_fa16(lay43_fa15_s, lay42_fa7_c, lay42_fa6_c, lay43_fa16_s, lay43_fa16_c);
wire lay43_fa17_s, lay43_fa17_c;
full_adder lay43_fa17(lay43_fa16_s, lay42_fa5_c, lay42_fa4_c, lay43_fa17_s, lay43_fa17_c);
wire lay43_fa18_s, lay43_fa18_c;
full_adder lay43_fa18(lay43_fa17_s, lay42_fa3_c, lay42_fa2_c, lay43_fa18_s, lay43_fa18_c);
wire lay43_fa19_s, lay43_fa19_c;
full_adder lay43_fa19(lay43_fa18_s, lay42_fa1_c, lay42_fa0_c, lay43_fa19_s, lay43_fa19_c);
assign prod[43] = lay43_fa19_s;

wire lay44_fa0_s, lay44_fa0_c;
full_adder lay44_fa0(a31b13, a30b14, a29b15, lay44_fa0_s, lay44_fa0_c);
wire lay44_fa1_s, lay44_fa1_c;
full_adder lay44_fa1(lay44_fa0_s, a28b16, a27b17, lay44_fa1_s, lay44_fa1_c);
wire lay44_fa2_s, lay44_fa2_c;
full_adder lay44_fa2(lay44_fa1_s, a26b18, a25b19, lay44_fa2_s, lay44_fa2_c);
wire lay44_fa3_s, lay44_fa3_c;
full_adder lay44_fa3(lay44_fa2_s, a24b20, a23b21, lay44_fa3_s, lay44_fa3_c);
wire lay44_fa4_s, lay44_fa4_c;
full_adder lay44_fa4(lay44_fa3_s, a22b22, a21b23, lay44_fa4_s, lay44_fa4_c);
wire lay44_fa5_s, lay44_fa5_c;
full_adder lay44_fa5(lay44_fa4_s, a20b24, a19b25, lay44_fa5_s, lay44_fa5_c);
wire lay44_fa6_s, lay44_fa6_c;
full_adder lay44_fa6(lay44_fa5_s, a18b26, a17b27, lay44_fa6_s, lay44_fa6_c);
wire lay44_fa7_s, lay44_fa7_c;
full_adder lay44_fa7(lay44_fa6_s, a16b28, a15b29, lay44_fa7_s, lay44_fa7_c);
wire lay44_fa8_s, lay44_fa8_c;
full_adder lay44_fa8(lay44_fa7_s, a14b30, a13b31, lay44_fa8_s, lay44_fa8_c);
wire lay44_fa9_s, lay44_fa9_c;
full_adder lay44_fa9(lay44_fa8_s, lay43_fa19_c, lay43_fa18_c, lay44_fa9_s, lay44_fa9_c);
wire lay44_fa10_s, lay44_fa10_c;
full_adder lay44_fa10(lay44_fa9_s, lay43_fa17_c, lay43_fa16_c, lay44_fa10_s, lay44_fa10_c);
wire lay44_fa11_s, lay44_fa11_c;
full_adder lay44_fa11(lay44_fa10_s, lay43_fa15_c, lay43_fa14_c, lay44_fa11_s, lay44_fa11_c);
wire lay44_fa12_s, lay44_fa12_c;
full_adder lay44_fa12(lay44_fa11_s, lay43_fa13_c, lay43_fa12_c, lay44_fa12_s, lay44_fa12_c);
wire lay44_fa13_s, lay44_fa13_c;
full_adder lay44_fa13(lay44_fa12_s, lay43_fa11_c, lay43_fa10_c, lay44_fa13_s, lay44_fa13_c);
wire lay44_fa14_s, lay44_fa14_c;
full_adder lay44_fa14(lay44_fa13_s, lay43_fa9_c, lay43_fa8_c, lay44_fa14_s, lay44_fa14_c);
wire lay44_fa15_s, lay44_fa15_c;
full_adder lay44_fa15(lay44_fa14_s, lay43_fa7_c, lay43_fa6_c, lay44_fa15_s, lay44_fa15_c);
wire lay44_fa16_s, lay44_fa16_c;
full_adder lay44_fa16(lay44_fa15_s, lay43_fa5_c, lay43_fa4_c, lay44_fa16_s, lay44_fa16_c);
wire lay44_fa17_s, lay44_fa17_c;
full_adder lay44_fa17(lay44_fa16_s, lay43_fa3_c, lay43_fa2_c, lay44_fa17_s, lay44_fa17_c);
wire lay44_fa18_s, lay44_fa18_c;
full_adder lay44_fa18(lay44_fa17_s, lay43_fa1_c, lay43_fa0_c, lay44_fa18_s, lay44_fa18_c);
assign prod[44] = lay44_fa18_s;

wire lay45_fa0_s, lay45_fa0_c;
full_adder lay45_fa0(a31b14, a30b15, a29b16, lay45_fa0_s, lay45_fa0_c);
wire lay45_fa1_s, lay45_fa1_c;
full_adder lay45_fa1(lay45_fa0_s, a28b17, a27b18, lay45_fa1_s, lay45_fa1_c);
wire lay45_fa2_s, lay45_fa2_c;
full_adder lay45_fa2(lay45_fa1_s, a26b19, a25b20, lay45_fa2_s, lay45_fa2_c);
wire lay45_fa3_s, lay45_fa3_c;
full_adder lay45_fa3(lay45_fa2_s, a24b21, a23b22, lay45_fa3_s, lay45_fa3_c);
wire lay45_fa4_s, lay45_fa4_c;
full_adder lay45_fa4(lay45_fa3_s, a22b23, a21b24, lay45_fa4_s, lay45_fa4_c);
wire lay45_fa5_s, lay45_fa5_c;
full_adder lay45_fa5(lay45_fa4_s, a20b25, a19b26, lay45_fa5_s, lay45_fa5_c);
wire lay45_fa6_s, lay45_fa6_c;
full_adder lay45_fa6(lay45_fa5_s, a18b27, a17b28, lay45_fa6_s, lay45_fa6_c);
wire lay45_fa7_s, lay45_fa7_c;
full_adder lay45_fa7(lay45_fa6_s, a16b29, a15b30, lay45_fa7_s, lay45_fa7_c);
wire lay45_fa8_s, lay45_fa8_c;
full_adder lay45_fa8(lay45_fa7_s, a14b31, lay44_fa18_c, lay45_fa8_s, lay45_fa8_c);
wire lay45_fa9_s, lay45_fa9_c;
full_adder lay45_fa9(lay45_fa8_s, lay44_fa17_c, lay44_fa16_c, lay45_fa9_s, lay45_fa9_c);
wire lay45_fa10_s, lay45_fa10_c;
full_adder lay45_fa10(lay45_fa9_s, lay44_fa15_c, lay44_fa14_c, lay45_fa10_s, lay45_fa10_c);
wire lay45_fa11_s, lay45_fa11_c;
full_adder lay45_fa11(lay45_fa10_s, lay44_fa13_c, lay44_fa12_c, lay45_fa11_s, lay45_fa11_c);
wire lay45_fa12_s, lay45_fa12_c;
full_adder lay45_fa12(lay45_fa11_s, lay44_fa11_c, lay44_fa10_c, lay45_fa12_s, lay45_fa12_c);
wire lay45_fa13_s, lay45_fa13_c;
full_adder lay45_fa13(lay45_fa12_s, lay44_fa9_c, lay44_fa8_c, lay45_fa13_s, lay45_fa13_c);
wire lay45_fa14_s, lay45_fa14_c;
full_adder lay45_fa14(lay45_fa13_s, lay44_fa7_c, lay44_fa6_c, lay45_fa14_s, lay45_fa14_c);
wire lay45_fa15_s, lay45_fa15_c;
full_adder lay45_fa15(lay45_fa14_s, lay44_fa5_c, lay44_fa4_c, lay45_fa15_s, lay45_fa15_c);
wire lay45_fa16_s, lay45_fa16_c;
full_adder lay45_fa16(lay45_fa15_s, lay44_fa3_c, lay44_fa2_c, lay45_fa16_s, lay45_fa16_c);
wire lay45_fa17_s, lay45_fa17_c;
full_adder lay45_fa17(lay45_fa16_s, lay44_fa1_c, lay44_fa0_c, lay45_fa17_s, lay45_fa17_c);
assign prod[45] = lay45_fa17_s;

wire lay46_fa0_s, lay46_fa0_c;
full_adder lay46_fa0(a31b15, a30b16, a29b17, lay46_fa0_s, lay46_fa0_c);
wire lay46_fa1_s, lay46_fa1_c;
full_adder lay46_fa1(lay46_fa0_s, a28b18, a27b19, lay46_fa1_s, lay46_fa1_c);
wire lay46_fa2_s, lay46_fa2_c;
full_adder lay46_fa2(lay46_fa1_s, a26b20, a25b21, lay46_fa2_s, lay46_fa2_c);
wire lay46_fa3_s, lay46_fa3_c;
full_adder lay46_fa3(lay46_fa2_s, a24b22, a23b23, lay46_fa3_s, lay46_fa3_c);
wire lay46_fa4_s, lay46_fa4_c;
full_adder lay46_fa4(lay46_fa3_s, a22b24, a21b25, lay46_fa4_s, lay46_fa4_c);
wire lay46_fa5_s, lay46_fa5_c;
full_adder lay46_fa5(lay46_fa4_s, a20b26, a19b27, lay46_fa5_s, lay46_fa5_c);
wire lay46_fa6_s, lay46_fa6_c;
full_adder lay46_fa6(lay46_fa5_s, a18b28, a17b29, lay46_fa6_s, lay46_fa6_c);
wire lay46_fa7_s, lay46_fa7_c;
full_adder lay46_fa7(lay46_fa6_s, a16b30, a15b31, lay46_fa7_s, lay46_fa7_c);
wire lay46_fa8_s, lay46_fa8_c;
full_adder lay46_fa8(lay46_fa7_s, lay45_fa17_c, lay45_fa16_c, lay46_fa8_s, lay46_fa8_c);
wire lay46_fa9_s, lay46_fa9_c;
full_adder lay46_fa9(lay46_fa8_s, lay45_fa15_c, lay45_fa14_c, lay46_fa9_s, lay46_fa9_c);
wire lay46_fa10_s, lay46_fa10_c;
full_adder lay46_fa10(lay46_fa9_s, lay45_fa13_c, lay45_fa12_c, lay46_fa10_s, lay46_fa10_c);
wire lay46_fa11_s, lay46_fa11_c;
full_adder lay46_fa11(lay46_fa10_s, lay45_fa11_c, lay45_fa10_c, lay46_fa11_s, lay46_fa11_c);
wire lay46_fa12_s, lay46_fa12_c;
full_adder lay46_fa12(lay46_fa11_s, lay45_fa9_c, lay45_fa8_c, lay46_fa12_s, lay46_fa12_c);
wire lay46_fa13_s, lay46_fa13_c;
full_adder lay46_fa13(lay46_fa12_s, lay45_fa7_c, lay45_fa6_c, lay46_fa13_s, lay46_fa13_c);
wire lay46_fa14_s, lay46_fa14_c;
full_adder lay46_fa14(lay46_fa13_s, lay45_fa5_c, lay45_fa4_c, lay46_fa14_s, lay46_fa14_c);
wire lay46_fa15_s, lay46_fa15_c;
full_adder lay46_fa15(lay46_fa14_s, lay45_fa3_c, lay45_fa2_c, lay46_fa15_s, lay46_fa15_c);
wire lay46_fa16_s, lay46_fa16_c;
full_adder lay46_fa16(lay46_fa15_s, lay45_fa1_c, lay45_fa0_c, lay46_fa16_s, lay46_fa16_c);
assign prod[46] = lay46_fa16_s;

wire lay47_fa0_s, lay47_fa0_c;
full_adder lay47_fa0(a31b16, a30b17, a29b18, lay47_fa0_s, lay47_fa0_c);
wire lay47_fa1_s, lay47_fa1_c;
full_adder lay47_fa1(lay47_fa0_s, a28b19, a27b20, lay47_fa1_s, lay47_fa1_c);
wire lay47_fa2_s, lay47_fa2_c;
full_adder lay47_fa2(lay47_fa1_s, a26b21, a25b22, lay47_fa2_s, lay47_fa2_c);
wire lay47_fa3_s, lay47_fa3_c;
full_adder lay47_fa3(lay47_fa2_s, a24b23, a23b24, lay47_fa3_s, lay47_fa3_c);
wire lay47_fa4_s, lay47_fa4_c;
full_adder lay47_fa4(lay47_fa3_s, a22b25, a21b26, lay47_fa4_s, lay47_fa4_c);
wire lay47_fa5_s, lay47_fa5_c;
full_adder lay47_fa5(lay47_fa4_s, a20b27, a19b28, lay47_fa5_s, lay47_fa5_c);
wire lay47_fa6_s, lay47_fa6_c;
full_adder lay47_fa6(lay47_fa5_s, a18b29, a17b30, lay47_fa6_s, lay47_fa6_c);
wire lay47_fa7_s, lay47_fa7_c;
full_adder lay47_fa7(lay47_fa6_s, a16b31, lay46_fa16_c, lay47_fa7_s, lay47_fa7_c);
wire lay47_fa8_s, lay47_fa8_c;
full_adder lay47_fa8(lay47_fa7_s, lay46_fa15_c, lay46_fa14_c, lay47_fa8_s, lay47_fa8_c);
wire lay47_fa9_s, lay47_fa9_c;
full_adder lay47_fa9(lay47_fa8_s, lay46_fa13_c, lay46_fa12_c, lay47_fa9_s, lay47_fa9_c);
wire lay47_fa10_s, lay47_fa10_c;
full_adder lay47_fa10(lay47_fa9_s, lay46_fa11_c, lay46_fa10_c, lay47_fa10_s, lay47_fa10_c);
wire lay47_fa11_s, lay47_fa11_c;
full_adder lay47_fa11(lay47_fa10_s, lay46_fa9_c, lay46_fa8_c, lay47_fa11_s, lay47_fa11_c);
wire lay47_fa12_s, lay47_fa12_c;
full_adder lay47_fa12(lay47_fa11_s, lay46_fa7_c, lay46_fa6_c, lay47_fa12_s, lay47_fa12_c);
wire lay47_fa13_s, lay47_fa13_c;
full_adder lay47_fa13(lay47_fa12_s, lay46_fa5_c, lay46_fa4_c, lay47_fa13_s, lay47_fa13_c);
wire lay47_fa14_s, lay47_fa14_c;
full_adder lay47_fa14(lay47_fa13_s, lay46_fa3_c, lay46_fa2_c, lay47_fa14_s, lay47_fa14_c);
wire lay47_fa15_s, lay47_fa15_c;
full_adder lay47_fa15(lay47_fa14_s, lay46_fa1_c, lay46_fa0_c, lay47_fa15_s, lay47_fa15_c);
assign prod[47] = lay47_fa15_s;

wire lay48_fa0_s, lay48_fa0_c;
full_adder lay48_fa0(a31b17, a30b18, a29b19, lay48_fa0_s, lay48_fa0_c);
wire lay48_fa1_s, lay48_fa1_c;
full_adder lay48_fa1(lay48_fa0_s, a28b20, a27b21, lay48_fa1_s, lay48_fa1_c);
wire lay48_fa2_s, lay48_fa2_c;
full_adder lay48_fa2(lay48_fa1_s, a26b22, a25b23, lay48_fa2_s, lay48_fa2_c);
wire lay48_fa3_s, lay48_fa3_c;
full_adder lay48_fa3(lay48_fa2_s, a24b24, a23b25, lay48_fa3_s, lay48_fa3_c);
wire lay48_fa4_s, lay48_fa4_c;
full_adder lay48_fa4(lay48_fa3_s, a22b26, a21b27, lay48_fa4_s, lay48_fa4_c);
wire lay48_fa5_s, lay48_fa5_c;
full_adder lay48_fa5(lay48_fa4_s, a20b28, a19b29, lay48_fa5_s, lay48_fa5_c);
wire lay48_fa6_s, lay48_fa6_c;
full_adder lay48_fa6(lay48_fa5_s, a18b30, a17b31, lay48_fa6_s, lay48_fa6_c);
wire lay48_fa7_s, lay48_fa7_c;
full_adder lay48_fa7(lay48_fa6_s, lay47_fa15_c, lay47_fa14_c, lay48_fa7_s, lay48_fa7_c);
wire lay48_fa8_s, lay48_fa8_c;
full_adder lay48_fa8(lay48_fa7_s, lay47_fa13_c, lay47_fa12_c, lay48_fa8_s, lay48_fa8_c);
wire lay48_fa9_s, lay48_fa9_c;
full_adder lay48_fa9(lay48_fa8_s, lay47_fa11_c, lay47_fa10_c, lay48_fa9_s, lay48_fa9_c);
wire lay48_fa10_s, lay48_fa10_c;
full_adder lay48_fa10(lay48_fa9_s, lay47_fa9_c, lay47_fa8_c, lay48_fa10_s, lay48_fa10_c);
wire lay48_fa11_s, lay48_fa11_c;
full_adder lay48_fa11(lay48_fa10_s, lay47_fa7_c, lay47_fa6_c, lay48_fa11_s, lay48_fa11_c);
wire lay48_fa12_s, lay48_fa12_c;
full_adder lay48_fa12(lay48_fa11_s, lay47_fa5_c, lay47_fa4_c, lay48_fa12_s, lay48_fa12_c);
wire lay48_fa13_s, lay48_fa13_c;
full_adder lay48_fa13(lay48_fa12_s, lay47_fa3_c, lay47_fa2_c, lay48_fa13_s, lay48_fa13_c);
wire lay48_fa14_s, lay48_fa14_c;
full_adder lay48_fa14(lay48_fa13_s, lay47_fa1_c, lay47_fa0_c, lay48_fa14_s, lay48_fa14_c);
assign prod[48] = lay48_fa14_s;

wire lay49_fa0_s, lay49_fa0_c;
full_adder lay49_fa0(a31b18, a30b19, a29b20, lay49_fa0_s, lay49_fa0_c);
wire lay49_fa1_s, lay49_fa1_c;
full_adder lay49_fa1(lay49_fa0_s, a28b21, a27b22, lay49_fa1_s, lay49_fa1_c);
wire lay49_fa2_s, lay49_fa2_c;
full_adder lay49_fa2(lay49_fa1_s, a26b23, a25b24, lay49_fa2_s, lay49_fa2_c);
wire lay49_fa3_s, lay49_fa3_c;
full_adder lay49_fa3(lay49_fa2_s, a24b25, a23b26, lay49_fa3_s, lay49_fa3_c);
wire lay49_fa4_s, lay49_fa4_c;
full_adder lay49_fa4(lay49_fa3_s, a22b27, a21b28, lay49_fa4_s, lay49_fa4_c);
wire lay49_fa5_s, lay49_fa5_c;
full_adder lay49_fa5(lay49_fa4_s, a20b29, a19b30, lay49_fa5_s, lay49_fa5_c);
wire lay49_fa6_s, lay49_fa6_c;
full_adder lay49_fa6(lay49_fa5_s, a18b31, lay48_fa14_c, lay49_fa6_s, lay49_fa6_c);
wire lay49_fa7_s, lay49_fa7_c;
full_adder lay49_fa7(lay49_fa6_s, lay48_fa13_c, lay48_fa12_c, lay49_fa7_s, lay49_fa7_c);
wire lay49_fa8_s, lay49_fa8_c;
full_adder lay49_fa8(lay49_fa7_s, lay48_fa11_c, lay48_fa10_c, lay49_fa8_s, lay49_fa8_c);
wire lay49_fa9_s, lay49_fa9_c;
full_adder lay49_fa9(lay49_fa8_s, lay48_fa9_c, lay48_fa8_c, lay49_fa9_s, lay49_fa9_c);
wire lay49_fa10_s, lay49_fa10_c;
full_adder lay49_fa10(lay49_fa9_s, lay48_fa7_c, lay48_fa6_c, lay49_fa10_s, lay49_fa10_c);
wire lay49_fa11_s, lay49_fa11_c;
full_adder lay49_fa11(lay49_fa10_s, lay48_fa5_c, lay48_fa4_c, lay49_fa11_s, lay49_fa11_c);
wire lay49_fa12_s, lay49_fa12_c;
full_adder lay49_fa12(lay49_fa11_s, lay48_fa3_c, lay48_fa2_c, lay49_fa12_s, lay49_fa12_c);
wire lay49_fa13_s, lay49_fa13_c;
full_adder lay49_fa13(lay49_fa12_s, lay48_fa1_c, lay48_fa0_c, lay49_fa13_s, lay49_fa13_c);
assign prod[49] = lay49_fa13_s;

wire lay50_fa0_s, lay50_fa0_c;
full_adder lay50_fa0(a31b19, a30b20, a29b21, lay50_fa0_s, lay50_fa0_c);
wire lay50_fa1_s, lay50_fa1_c;
full_adder lay50_fa1(lay50_fa0_s, a28b22, a27b23, lay50_fa1_s, lay50_fa1_c);
wire lay50_fa2_s, lay50_fa2_c;
full_adder lay50_fa2(lay50_fa1_s, a26b24, a25b25, lay50_fa2_s, lay50_fa2_c);
wire lay50_fa3_s, lay50_fa3_c;
full_adder lay50_fa3(lay50_fa2_s, a24b26, a23b27, lay50_fa3_s, lay50_fa3_c);
wire lay50_fa4_s, lay50_fa4_c;
full_adder lay50_fa4(lay50_fa3_s, a22b28, a21b29, lay50_fa4_s, lay50_fa4_c);
wire lay50_fa5_s, lay50_fa5_c;
full_adder lay50_fa5(lay50_fa4_s, a20b30, a19b31, lay50_fa5_s, lay50_fa5_c);
wire lay50_fa6_s, lay50_fa6_c;
full_adder lay50_fa6(lay50_fa5_s, lay49_fa13_c, lay49_fa12_c, lay50_fa6_s, lay50_fa6_c);
wire lay50_fa7_s, lay50_fa7_c;
full_adder lay50_fa7(lay50_fa6_s, lay49_fa11_c, lay49_fa10_c, lay50_fa7_s, lay50_fa7_c);
wire lay50_fa8_s, lay50_fa8_c;
full_adder lay50_fa8(lay50_fa7_s, lay49_fa9_c, lay49_fa8_c, lay50_fa8_s, lay50_fa8_c);
wire lay50_fa9_s, lay50_fa9_c;
full_adder lay50_fa9(lay50_fa8_s, lay49_fa7_c, lay49_fa6_c, lay50_fa9_s, lay50_fa9_c);
wire lay50_fa10_s, lay50_fa10_c;
full_adder lay50_fa10(lay50_fa9_s, lay49_fa5_c, lay49_fa4_c, lay50_fa10_s, lay50_fa10_c);
wire lay50_fa11_s, lay50_fa11_c;
full_adder lay50_fa11(lay50_fa10_s, lay49_fa3_c, lay49_fa2_c, lay50_fa11_s, lay50_fa11_c);
wire lay50_fa12_s, lay50_fa12_c;
full_adder lay50_fa12(lay50_fa11_s, lay49_fa1_c, lay49_fa0_c, lay50_fa12_s, lay50_fa12_c);
assign prod[50] = lay50_fa12_s;

wire lay51_fa0_s, lay51_fa0_c;
full_adder lay51_fa0(a31b20, a30b21, a29b22, lay51_fa0_s, lay51_fa0_c);
wire lay51_fa1_s, lay51_fa1_c;
full_adder lay51_fa1(lay51_fa0_s, a28b23, a27b24, lay51_fa1_s, lay51_fa1_c);
wire lay51_fa2_s, lay51_fa2_c;
full_adder lay51_fa2(lay51_fa1_s, a26b25, a25b26, lay51_fa2_s, lay51_fa2_c);
wire lay51_fa3_s, lay51_fa3_c;
full_adder lay51_fa3(lay51_fa2_s, a24b27, a23b28, lay51_fa3_s, lay51_fa3_c);
wire lay51_fa4_s, lay51_fa4_c;
full_adder lay51_fa4(lay51_fa3_s, a22b29, a21b30, lay51_fa4_s, lay51_fa4_c);
wire lay51_fa5_s, lay51_fa5_c;
full_adder lay51_fa5(lay51_fa4_s, a20b31, lay50_fa12_c, lay51_fa5_s, lay51_fa5_c);
wire lay51_fa6_s, lay51_fa6_c;
full_adder lay51_fa6(lay51_fa5_s, lay50_fa11_c, lay50_fa10_c, lay51_fa6_s, lay51_fa6_c);
wire lay51_fa7_s, lay51_fa7_c;
full_adder lay51_fa7(lay51_fa6_s, lay50_fa9_c, lay50_fa8_c, lay51_fa7_s, lay51_fa7_c);
wire lay51_fa8_s, lay51_fa8_c;
full_adder lay51_fa8(lay51_fa7_s, lay50_fa7_c, lay50_fa6_c, lay51_fa8_s, lay51_fa8_c);
wire lay51_fa9_s, lay51_fa9_c;
full_adder lay51_fa9(lay51_fa8_s, lay50_fa5_c, lay50_fa4_c, lay51_fa9_s, lay51_fa9_c);
wire lay51_fa10_s, lay51_fa10_c;
full_adder lay51_fa10(lay51_fa9_s, lay50_fa3_c, lay50_fa2_c, lay51_fa10_s, lay51_fa10_c);
wire lay51_fa11_s, lay51_fa11_c;
full_adder lay51_fa11(lay51_fa10_s, lay50_fa1_c, lay50_fa0_c, lay51_fa11_s, lay51_fa11_c);
assign prod[51] = lay51_fa11_s;

wire lay52_fa0_s, lay52_fa0_c;
full_adder lay52_fa0(a31b21, a30b22, a29b23, lay52_fa0_s, lay52_fa0_c);
wire lay52_fa1_s, lay52_fa1_c;
full_adder lay52_fa1(lay52_fa0_s, a28b24, a27b25, lay52_fa1_s, lay52_fa1_c);
wire lay52_fa2_s, lay52_fa2_c;
full_adder lay52_fa2(lay52_fa1_s, a26b26, a25b27, lay52_fa2_s, lay52_fa2_c);
wire lay52_fa3_s, lay52_fa3_c;
full_adder lay52_fa3(lay52_fa2_s, a24b28, a23b29, lay52_fa3_s, lay52_fa3_c);
wire lay52_fa4_s, lay52_fa4_c;
full_adder lay52_fa4(lay52_fa3_s, a22b30, a21b31, lay52_fa4_s, lay52_fa4_c);
wire lay52_fa5_s, lay52_fa5_c;
full_adder lay52_fa5(lay52_fa4_s, lay51_fa11_c, lay51_fa10_c, lay52_fa5_s, lay52_fa5_c);
wire lay52_fa6_s, lay52_fa6_c;
full_adder lay52_fa6(lay52_fa5_s, lay51_fa9_c, lay51_fa8_c, lay52_fa6_s, lay52_fa6_c);
wire lay52_fa7_s, lay52_fa7_c;
full_adder lay52_fa7(lay52_fa6_s, lay51_fa7_c, lay51_fa6_c, lay52_fa7_s, lay52_fa7_c);
wire lay52_fa8_s, lay52_fa8_c;
full_adder lay52_fa8(lay52_fa7_s, lay51_fa5_c, lay51_fa4_c, lay52_fa8_s, lay52_fa8_c);
wire lay52_fa9_s, lay52_fa9_c;
full_adder lay52_fa9(lay52_fa8_s, lay51_fa3_c, lay51_fa2_c, lay52_fa9_s, lay52_fa9_c);
wire lay52_fa10_s, lay52_fa10_c;
full_adder lay52_fa10(lay52_fa9_s, lay51_fa1_c, lay51_fa0_c, lay52_fa10_s, lay52_fa10_c);
assign prod[52] = lay52_fa10_s;

wire lay53_fa0_s, lay53_fa0_c;
full_adder lay53_fa0(a31b22, a30b23, a29b24, lay53_fa0_s, lay53_fa0_c);
wire lay53_fa1_s, lay53_fa1_c;
full_adder lay53_fa1(lay53_fa0_s, a28b25, a27b26, lay53_fa1_s, lay53_fa1_c);
wire lay53_fa2_s, lay53_fa2_c;
full_adder lay53_fa2(lay53_fa1_s, a26b27, a25b28, lay53_fa2_s, lay53_fa2_c);
wire lay53_fa3_s, lay53_fa3_c;
full_adder lay53_fa3(lay53_fa2_s, a24b29, a23b30, lay53_fa3_s, lay53_fa3_c);
wire lay53_fa4_s, lay53_fa4_c;
full_adder lay53_fa4(lay53_fa3_s, a22b31, lay52_fa10_c, lay53_fa4_s, lay53_fa4_c);
wire lay53_fa5_s, lay53_fa5_c;
full_adder lay53_fa5(lay53_fa4_s, lay52_fa9_c, lay52_fa8_c, lay53_fa5_s, lay53_fa5_c);
wire lay53_fa6_s, lay53_fa6_c;
full_adder lay53_fa6(lay53_fa5_s, lay52_fa7_c, lay52_fa6_c, lay53_fa6_s, lay53_fa6_c);
wire lay53_fa7_s, lay53_fa7_c;
full_adder lay53_fa7(lay53_fa6_s, lay52_fa5_c, lay52_fa4_c, lay53_fa7_s, lay53_fa7_c);
wire lay53_fa8_s, lay53_fa8_c;
full_adder lay53_fa8(lay53_fa7_s, lay52_fa3_c, lay52_fa2_c, lay53_fa8_s, lay53_fa8_c);
wire lay53_fa9_s, lay53_fa9_c;
full_adder lay53_fa9(lay53_fa8_s, lay52_fa1_c, lay52_fa0_c, lay53_fa9_s, lay53_fa9_c);
assign prod[53] = lay53_fa9_s;

wire lay54_fa0_s, lay54_fa0_c;
full_adder lay54_fa0(a31b23, a30b24, a29b25, lay54_fa0_s, lay54_fa0_c);
wire lay54_fa1_s, lay54_fa1_c;
full_adder lay54_fa1(lay54_fa0_s, a28b26, a27b27, lay54_fa1_s, lay54_fa1_c);
wire lay54_fa2_s, lay54_fa2_c;
full_adder lay54_fa2(lay54_fa1_s, a26b28, a25b29, lay54_fa2_s, lay54_fa2_c);
wire lay54_fa3_s, lay54_fa3_c;
full_adder lay54_fa3(lay54_fa2_s, a24b30, a23b31, lay54_fa3_s, lay54_fa3_c);
wire lay54_fa4_s, lay54_fa4_c;
full_adder lay54_fa4(lay54_fa3_s, lay53_fa9_c, lay53_fa8_c, lay54_fa4_s, lay54_fa4_c);
wire lay54_fa5_s, lay54_fa5_c;
full_adder lay54_fa5(lay54_fa4_s, lay53_fa7_c, lay53_fa6_c, lay54_fa5_s, lay54_fa5_c);
wire lay54_fa6_s, lay54_fa6_c;
full_adder lay54_fa6(lay54_fa5_s, lay53_fa5_c, lay53_fa4_c, lay54_fa6_s, lay54_fa6_c);
wire lay54_fa7_s, lay54_fa7_c;
full_adder lay54_fa7(lay54_fa6_s, lay53_fa3_c, lay53_fa2_c, lay54_fa7_s, lay54_fa7_c);
wire lay54_fa8_s, lay54_fa8_c;
full_adder lay54_fa8(lay54_fa7_s, lay53_fa1_c, lay53_fa0_c, lay54_fa8_s, lay54_fa8_c);
assign prod[54] = lay54_fa8_s;

wire lay55_fa0_s, lay55_fa0_c;
full_adder lay55_fa0(a31b24, a30b25, a29b26, lay55_fa0_s, lay55_fa0_c);
wire lay55_fa1_s, lay55_fa1_c;
full_adder lay55_fa1(lay55_fa0_s, a28b27, a27b28, lay55_fa1_s, lay55_fa1_c);
wire lay55_fa2_s, lay55_fa2_c;
full_adder lay55_fa2(lay55_fa1_s, a26b29, a25b30, lay55_fa2_s, lay55_fa2_c);
wire lay55_fa3_s, lay55_fa3_c;
full_adder lay55_fa3(lay55_fa2_s, a24b31, lay54_fa8_c, lay55_fa3_s, lay55_fa3_c);
wire lay55_fa4_s, lay55_fa4_c;
full_adder lay55_fa4(lay55_fa3_s, lay54_fa7_c, lay54_fa6_c, lay55_fa4_s, lay55_fa4_c);
wire lay55_fa5_s, lay55_fa5_c;
full_adder lay55_fa5(lay55_fa4_s, lay54_fa5_c, lay54_fa4_c, lay55_fa5_s, lay55_fa5_c);
wire lay55_fa6_s, lay55_fa6_c;
full_adder lay55_fa6(lay55_fa5_s, lay54_fa3_c, lay54_fa2_c, lay55_fa6_s, lay55_fa6_c);
wire lay55_fa7_s, lay55_fa7_c;
full_adder lay55_fa7(lay55_fa6_s, lay54_fa1_c, lay54_fa0_c, lay55_fa7_s, lay55_fa7_c);
assign prod[55] = lay55_fa7_s;

wire lay56_fa0_s, lay56_fa0_c;
full_adder lay56_fa0(a31b25, a30b26, a29b27, lay56_fa0_s, lay56_fa0_c);
wire lay56_fa1_s, lay56_fa1_c;
full_adder lay56_fa1(lay56_fa0_s, a28b28, a27b29, lay56_fa1_s, lay56_fa1_c);
wire lay56_fa2_s, lay56_fa2_c;
full_adder lay56_fa2(lay56_fa1_s, a26b30, a25b31, lay56_fa2_s, lay56_fa2_c);
wire lay56_fa3_s, lay56_fa3_c;
full_adder lay56_fa3(lay56_fa2_s, lay55_fa7_c, lay55_fa6_c, lay56_fa3_s, lay56_fa3_c);
wire lay56_fa4_s, lay56_fa4_c;
full_adder lay56_fa4(lay56_fa3_s, lay55_fa5_c, lay55_fa4_c, lay56_fa4_s, lay56_fa4_c);
wire lay56_fa5_s, lay56_fa5_c;
full_adder lay56_fa5(lay56_fa4_s, lay55_fa3_c, lay55_fa2_c, lay56_fa5_s, lay56_fa5_c);
wire lay56_fa6_s, lay56_fa6_c;
full_adder lay56_fa6(lay56_fa5_s, lay55_fa1_c, lay55_fa0_c, lay56_fa6_s, lay56_fa6_c);
assign prod[56] = lay56_fa6_s;

wire lay57_fa0_s, lay57_fa0_c;
full_adder lay57_fa0(a31b26, a30b27, a29b28, lay57_fa0_s, lay57_fa0_c);
wire lay57_fa1_s, lay57_fa1_c;
full_adder lay57_fa1(lay57_fa0_s, a28b29, a27b30, lay57_fa1_s, lay57_fa1_c);
wire lay57_fa2_s, lay57_fa2_c;
full_adder lay57_fa2(lay57_fa1_s, a26b31, lay56_fa6_c, lay57_fa2_s, lay57_fa2_c);
wire lay57_fa3_s, lay57_fa3_c;
full_adder lay57_fa3(lay57_fa2_s, lay56_fa5_c, lay56_fa4_c, lay57_fa3_s, lay57_fa3_c);
wire lay57_fa4_s, lay57_fa4_c;
full_adder lay57_fa4(lay57_fa3_s, lay56_fa3_c, lay56_fa2_c, lay57_fa4_s, lay57_fa4_c);
wire lay57_fa5_s, lay57_fa5_c;
full_adder lay57_fa5(lay57_fa4_s, lay56_fa1_c, lay56_fa0_c, lay57_fa5_s, lay57_fa5_c);
assign prod[57] = lay57_fa5_s;

wire lay58_fa0_s, lay58_fa0_c;
full_adder lay58_fa0(a31b27, a30b28, a29b29, lay58_fa0_s, lay58_fa0_c);
wire lay58_fa1_s, lay58_fa1_c;
full_adder lay58_fa1(lay58_fa0_s, a28b30, a27b31, lay58_fa1_s, lay58_fa1_c);
wire lay58_fa2_s, lay58_fa2_c;
full_adder lay58_fa2(lay58_fa1_s, lay57_fa5_c, lay57_fa4_c, lay58_fa2_s, lay58_fa2_c);
wire lay58_fa3_s, lay58_fa3_c;
full_adder lay58_fa3(lay58_fa2_s, lay57_fa3_c, lay57_fa2_c, lay58_fa3_s, lay58_fa3_c);
wire lay58_fa4_s, lay58_fa4_c;
full_adder lay58_fa4(lay58_fa3_s, lay57_fa1_c, lay57_fa0_c, lay58_fa4_s, lay58_fa4_c);
assign prod[58] = lay58_fa4_s;

wire lay59_fa0_s, lay59_fa0_c;
full_adder lay59_fa0(a31b28, a30b29, a29b30, lay59_fa0_s, lay59_fa0_c);
wire lay59_fa1_s, lay59_fa1_c;
full_adder lay59_fa1(lay59_fa0_s, a28b31, lay58_fa4_c, lay59_fa1_s, lay59_fa1_c);
wire lay59_fa2_s, lay59_fa2_c;
full_adder lay59_fa2(lay59_fa1_s, lay58_fa3_c, lay58_fa2_c, lay59_fa2_s, lay59_fa2_c);
wire lay59_fa3_s, lay59_fa3_c;
full_adder lay59_fa3(lay59_fa2_s, lay58_fa1_c, lay58_fa0_c, lay59_fa3_s, lay59_fa3_c);
assign prod[59] = lay59_fa3_s;

wire lay60_fa0_s, lay60_fa0_c;
full_adder lay60_fa0(a31b29, a30b30, a29b31, lay60_fa0_s, lay60_fa0_c);
wire lay60_fa1_s, lay60_fa1_c;
full_adder lay60_fa1(lay60_fa0_s, lay59_fa3_c, lay59_fa2_c, lay60_fa1_s, lay60_fa1_c);
wire lay60_fa2_s, lay60_fa2_c;
full_adder lay60_fa2(lay60_fa1_s, lay59_fa1_c, lay59_fa0_c, lay60_fa2_s, lay60_fa2_c);
assign prod[60] = lay60_fa2_s;

wire lay61_fa0_s, lay61_fa0_c;
full_adder lay61_fa0(a31b30, a30b31, lay60_fa2_c, lay61_fa0_s, lay61_fa0_c);
wire lay61_fa1_s, lay61_fa1_c;
full_adder lay61_fa1(lay61_fa0_s, lay60_fa1_c, lay60_fa0_c, lay61_fa1_s, lay61_fa1_c);
assign prod[61] = lay61_fa1_s;

wire lay62_fa0_s, lay62_fa0_c;
full_adder lay62_fa0(a31b31, lay61_fa1_c, lay61_fa0_c, lay62_fa0_s, lay62_fa0_c);
assign prod[62] = lay62_fa0_s;

wire lay63_ha0_s, lay63_ha0_c;
half_adder lay63_ha0(1'b1, lay62_fa0_c, lay63_ha0_s, lay63_ha0_c);
assign prod[63] = lay63_ha0_s;

//assign prod[63] = lay63_ha0_c;
assign prod_trim[31:0] = prod[31:0];


wire chk, chka, chkb, chkneg, chkpos;


//1 if all 1's
and neg_and(chkneg, prod[32], prod[33], prod[34], prod[35], prod[36], prod[37], prod[38], prod[39], prod[40], prod[41], prod[42], prod[43], prod[44], prod[45], prod[46], prod[47], prod[48], prod[49], prod[50], prod[51], prod[52], prod[53], prod[54], prod[55], prod[56], prod[57], prod[58], prod[59], prod[60], prod[61], prod[62], prod[63]);

//1 if all 0's 
nor pos_nor(chkpos, prod[32], prod[33], prod[34], prod[35], prod[36], prod[37], prod[38], prod[39], prod[40], prod[41], prod[42], prod[43], prod[44], prod[45], prod[46], prod[47], prod[48], prod[49], prod[50], prod[51], prod[52], prod[53], prod[54], prod[55], prod[56], prod[57], prod[58], prod[59], prod[60], prod[61], prod[62], prod[63]);

//1 if 0, 0 if nonzero
nor exc_check(chk, prod[0], prod[1], prod[2], prod[3], prod[4], prod[5], prod[6], prod[7], prod[8], prod[9], prod[10], prod[11], prod[12], prod[13], prod[14], prod[15], prod[16], prod[17], prod[18], prod[19], prod[20], prod[21], prod[22], prod[23], prod[24], prod[25], prod[26], prod[27], prod[28], prod[29], prod[30], prod[31]);

nor a_check(chka, a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17], a[18], a[19], a[20], a[21], a[22], a[23], a[24], a[25], a[26], a[27], a[28], a[29], a[30], a[31]);

nor b_check(chkb, b[0], b[1], b[2], b[3], b[4], b[5], b[6], b[7], b[8], b[9], b[10], b[11], b[12], b[13], b[14], b[15], b[16], b[17], b[18], b[19], b[20], b[21], b[22], b[23], b[24], b[25], b[26], b[27], b[28], b[29], b[30], b[31]);

wire non_zero, not_same, no_ovf;
//or ab_chk(non_zero, a_check, b_check)'

and exc(non_zero, chk, !chka, !chkb);

xnor ovf_and(no_ovf, chkneg, chkpos);

xor sign_xor(not_same, prod[63], prod_trim[31]);

or throw(exp, non_zero, not_same, no_ovf); 



endmodule