module lshift_1(A, out);
    input [31:0] A;
    output [31:0] out;

    assign out[0] = 0;
    assign out[1] = A[0];
    assign out[2] = A[1];
    assign out[3] = A[2];
    assign out[4] = A[3];
    assign out[5] = A[4];
    assign out[6] = A[5];
    assign out[7] = A[6];
    assign out[8] = A[7];
    assign out[9] = A[8];
    assign out[10] = A[9];
    assign out[11] = A[10];
    assign out[12] = A[11];
    assign out[13] = A[12];
    assign out[14] = A[13];
    assign out[15] = A[14];
    assign out[16] = A[15];
    assign out[17] = A[16];
    assign out[18] = A[17];
    assign out[19] = A[18];
    assign out[20] = A[19];
    assign out[21] = A[20];
    assign out[22] = A[21];
    assign out[23] = A[22];
    assign out[24] = A[23];
    assign out[25] = A[24];
    assign out[26] = A[25];
    assign out[27] = A[26];
    assign out[28] = A[27];
    assign out[29] = A[28];
    assign out[30] = A[29];
    assign out[31] = A[30];

endmodule


module lshift_2(A, out);
    input [31:0] A;
    output [31:0] out;


    assign out[0] = 0;
    assign out[1] = 0;
    assign out[2] = A[0];
    assign out[3] = A[1];
    assign out[4] = A[2];
    assign out[5] = A[3];
    assign out[6] = A[4];
    assign out[7] = A[5];
    assign out[8] = A[6];
    assign out[9] = A[7];
    assign out[10] = A[8];
    assign out[11] = A[9];
    assign out[12] = A[10];
    assign out[13] = A[11];
    assign out[14] = A[12];
    assign out[15] = A[13];
    assign out[16] = A[14];
    assign out[17] = A[15];
    assign out[18] = A[16];
    assign out[19] = A[17];
    assign out[20] = A[18];
    assign out[21] = A[19];
    assign out[22] = A[20];
    assign out[23] = A[21];
    assign out[24] = A[22];
    assign out[25] = A[23];
    assign out[26] = A[24];
    assign out[27] = A[25];
    assign out[28] = A[26];
    assign out[29] = A[27];
    assign out[30] = A[28];
    assign out[31] = A[29];

endmodule

module  lshift_4(A, out);
    input [31:0] A;
    output [31:0] out;


    assign out[0] = 0;
    assign out[1] = 0;
    assign out[2] = 0;
    assign out[3] = 0;
    assign out[4] = A[0];
    assign out[5] = A[1];
    assign out[6] = A[2];
    assign out[7] = A[3];
    assign out[8] = A[4];
    assign out[9] = A[5];
    assign out[10] = A[6];
    assign out[11] = A[7];
    assign out[12] = A[8];
    assign out[13] = A[9];
    assign out[14] = A[10];
    assign out[15] = A[11];
    assign out[16] = A[12];
    assign out[17] = A[13];
    assign out[18] = A[14];
    assign out[19] = A[15];
    assign out[20] = A[16];
    assign out[21] = A[17];
    assign out[22] = A[18];
    assign out[23] = A[19];
    assign out[24] = A[20];
    assign out[25] = A[21];
    assign out[26] = A[22];
    assign out[27] = A[23];
    assign out[28] = A[24];
    assign out[29] = A[25];
    assign out[30] = A[26];
    assign out[31] = A[27];

endmodule

module  lshift_8(A, out);
    input [31:0] A;
    output [31:0] out;

    assign out[0] = 0;
    assign out[1] = 0;
    assign out[2] = 0;
    assign out[3] = 0;
    assign out[4] = 0;
    assign out[5] = 0;
    assign out[6] = 0;
    assign out[7] = 0;
    assign out[8] = A[0];
    assign out[9] = A[1];
    assign out[10] = A[2];
    assign out[11] = A[3];
    assign out[12] = A[4];
    assign out[13] = A[5];
    assign out[14] = A[6];
    assign out[15] = A[7];
    assign out[16] = A[8];
    assign out[17] = A[9];
    assign out[18] = A[10];
    assign out[19] = A[11];
    assign out[20] = A[12];
    assign out[21] = A[13];
    assign out[22] = A[14];
    assign out[23] = A[15];
    assign out[24] = A[16];
    assign out[25] = A[17];
    assign out[26] = A[18];
    assign out[27] = A[19];
    assign out[28] = A[20];
    assign out[29] = A[21];
    assign out[30] = A[22];
    assign out[31] = A[23];

endmodule

module  lshift_16(A, out);
    input [31:0] A;
    output [31:0] out;

    assign out[0] = 0;
    assign out[1] = 0;
    assign out[2] = 0;
    assign out[3] = 0;
    assign out[4] = 0;
    assign out[5] = 0;
    assign out[6] = 0;
    assign out[7] = 0;
    assign out[8] = 0;
    assign out[9] = 0;
    assign out[10] = 0;
    assign out[11] = 0;
    assign out[12] = 0;
    assign out[13] = 0;
    assign out[14] = 0;
    assign out[15] = 0;
    assign out[16] = A[0];
    assign out[17] = A[1];
    assign out[18] = A[2];
    assign out[19] = A[3];
    assign out[20] = A[4];
    assign out[21] = A[5];
    assign out[22] = A[6];
    assign out[23] = A[7];
    assign out[24] = A[8];
    assign out[25] = A[9];
    assign out[26] = A[10];
    assign out[27] = A[11];
    assign out[28] = A[12];
    assign out[29] = A[13];
    assign out[30] = A[14];
    assign out[31] = A[15];

endmodule

module lshifter (A, shift_amt, out);
    input [31:0] A;
    input [4:0] shift_amt;

    output [31:0] out;
    wire [31:0] out_16, out_8, out_4, out_2, out_1, out_temp_1, out_temp_2, out_temp_3, out_temp_4;


    lshift_16 lshift_16(A, out_16);
    mux_2 mux_2_0(out_temp_1, shift_amt[4], A, out_16);
    lshift_8 lshift_8(out_temp_1, out_8);
    mux_2 mux_2_1(out_temp_2, shift_amt[3], out_temp_1, out_8);
    lshift_4 lshift_4(out_temp_2, out_4);
    mux_2 mux_2_2(out_temp_3, shift_amt[2], out_temp_2, out_4);
    lshift_2 lshift_2(out_temp_3, out_2);
    mux_2 mux_2_3(out_temp_4, shift_amt[1], out_temp_3, out_2);
    lshift_1 lshift_1(out_temp_4, out_1);
    mux_2 mux_2_4(out, shift_amt[0], out_temp_4, out_1);


endmodule