module rshift_1(A, out);
    input [31:0] A;
    output [31:0] out;

    assign out[0] = A[1];
    assign out[1] = A[2];
    assign out[2] = A[3];
    assign out[3] = A[4];
    assign out[4] = A[5];
    assign out[5] = A[6];
    assign out[6] = A[7];
    assign out[7] = A[8];
    assign out[8] = A[9];
    assign out[9] = A[10];
    assign out[10] = A[11];
    assign out[11] = A[12];
    assign out[12] = A[13];
    assign out[13] = A[14];
    assign out[14] = A[15];
    assign out[15] = A[16];
    assign out[16] = A[17];
    assign out[17] = A[18];
    assign out[18] = A[19];
    assign out[19] = A[20];
    assign out[20] = A[21];
    assign out[21] = A[22];
    assign out[22] = A[23];
    assign out[23] = A[24];
    assign out[24] = A[25];
    assign out[25] = A[26];
    assign out[26] = A[27];
    assign out[27] = A[28];
    assign out[28] = A[29];
    assign out[29] = A[30];
    assign out[30] = A[31];
    assign out[31] = A[31];

endmodule


module rshift_2(A, out);
    input [31:0] A;
    output [31:0] out;

    assign out[0] = A[2];
    assign out[1] = A[3];
    assign out[2] = A[4];
    assign out[3] = A[5];
    assign out[4] = A[6];
    assign out[5] = A[7];
    assign out[6] = A[8];
    assign out[7] = A[9];
    assign out[8] = A[10];
    assign out[9] = A[11];
    assign out[10] = A[12];
    assign out[11] = A[13];
    assign out[12] = A[14];
    assign out[13] = A[15];
    assign out[14] = A[16];
    assign out[15] = A[17];
    assign out[16] = A[18];
    assign out[17] = A[19];
    assign out[18] = A[20];
    assign out[19] = A[21];
    assign out[20] = A[22];
    assign out[21] = A[23];
    assign out[22] = A[24];
    assign out[23] = A[25];
    assign out[24] = A[26];
    assign out[25] = A[27];
    assign out[26] = A[28];
    assign out[27] = A[29];
    assign out[28] = A[30];
    assign out[29] = A[31];
    assign out[30] = A[31];
    assign out[31] = A[31];

endmodule

module  rshift_4(A, out);
    input [31:0] A;
    output [31:0] out;

    assign out[0] = A[4];
    assign out[1] = A[5];
    assign out[2] = A[6];
    assign out[3] = A[7];
    assign out[4] = A[8];
    assign out[5] = A[9];
    assign out[6] = A[10];
    assign out[7] = A[11];
    assign out[8] = A[12];
    assign out[9] = A[13];
    assign out[10] = A[14];
    assign out[11] = A[15];
    assign out[12] = A[16];
    assign out[13] = A[17];
    assign out[14] = A[18];
    assign out[15] = A[19];
    assign out[16] = A[20];
    assign out[17] = A[21];
    assign out[18] = A[22];
    assign out[19] = A[23];
    assign out[20] = A[24];
    assign out[21] = A[25];
    assign out[22] = A[26];
    assign out[23] = A[27];
    assign out[24] = A[28];
    assign out[25] = A[29];
    assign out[26] = A[30];
    assign out[27] = A[31];
    assign out[28] = A[31];
    assign out[29] = A[31];
    assign out[30] = A[31];
    assign out[31] = A[31];

endmodule

module  rshift_8(A, out);
    input [31:0] A;
    output [31:0] out;

    assign out[0] = A[8];
    assign out[1] = A[9];
    assign out[2] = A[10];
    assign out[3] = A[11];
    assign out[4] = A[12];
    assign out[5] = A[13];
    assign out[6] = A[14];
    assign out[7] = A[15];
    assign out[8] = A[16];
    assign out[9] = A[17];
    assign out[10] = A[18];
    assign out[11] = A[19];
    assign out[12] = A[20];
    assign out[13] = A[21];
    assign out[14] = A[22];
    assign out[15] = A[23];
    assign out[16] = A[24];
    assign out[17] = A[25];
    assign out[18] = A[26];
    assign out[19] = A[27];
    assign out[20] = A[28];
    assign out[21] = A[29];
    assign out[22] = A[30];
    assign out[23] = A[31];
    assign out[24] = A[31];
    assign out[25] = A[31];
    assign out[26] = A[31];
    assign out[27] = A[31];
    assign out[28] = A[31];
    assign out[29] = A[31];
    assign out[30] = A[31];
    assign out[31] = A[31];

endmodule

module  rshift_16(A, out);
    input [31:0] A;
    output [31:0] out;

    assign out[0] = A[16];
    assign out[1] = A[17];
    assign out[2] = A[18];
    assign out[3] = A[19];
    assign out[4] = A[20];
    assign out[5] = A[21];
    assign out[6] = A[22];
    assign out[7] = A[23];
    assign out[8] = A[24];
    assign out[9] = A[25];
    assign out[10] = A[26];
    assign out[11] = A[27];
    assign out[12] = A[28];
    assign out[13] = A[29];
    assign out[14] = A[30];
    assign out[15] = A[31];
    assign out[16] = A[31];
    assign out[17] = A[31];
    assign out[18] = A[31];
    assign out[19] = A[31];
    assign out[20] = A[31];
    assign out[21] = A[31];
    assign out[22] = A[31];
    assign out[23] = A[31];
    assign out[24] = A[31];
    assign out[25] = A[31];
    assign out[26] = A[31];
    assign out[27] = A[31];
    assign out[28] = A[31];
    assign out[29] = A[31];
    assign out[30] = A[31];
    assign out[31] = A[31];

endmodule

module rshifter (A, shift_amt, out);
    input [31:0] A;
    input [4:0] shift_amt;

    output [31:0] out;
    wire [31:0] out_16, out_8, out_4, out_2, out_1, out_temp_1, out_temp_2, out_temp_3, out_temp_4;


    rshift_16 rshift_16(A, out_16);
    mux_2 mux_2_0(out_temp_1, shift_amt[4], A, out_16);
    rshift_8 rshift_8(out_temp_1, out_8);
    mux_2 mux_2_1(out_temp_2, shift_amt[3], out_temp_1, out_8);
    rshift_4 rshift_4(out_temp_2, out_4);
    mux_2 mux_2_2(out_temp_3, shift_amt[2], out_temp_2, out_4);
    rshift_2 rshift_2(out_temp_3, out_2);
    mux_2 mux_2_3(out_temp_4, shift_amt[1], out_temp_3, out_2);
    rshift_1 rshift_1(out_temp_4, out_1);
    mux_2 mux_2_4(out, shift_amt[0], out_temp_4, out_1);


endmodule